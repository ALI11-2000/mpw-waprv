magic
tech sky130B
magscale 1 2
timestamp 1662898439
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2128 98808 97424
<< metal2 >>
rect 1398 99200 1454 100000
rect 3422 99200 3478 100000
rect 5446 99200 5502 100000
rect 7470 99200 7526 100000
rect 9494 99200 9550 100000
rect 11518 99200 11574 100000
rect 13542 99200 13598 100000
rect 15566 99200 15622 100000
rect 17590 99200 17646 100000
rect 19614 99200 19670 100000
rect 21638 99200 21694 100000
rect 23662 99200 23718 100000
rect 25686 99200 25742 100000
rect 27710 99200 27766 100000
rect 29734 99200 29790 100000
rect 31758 99200 31814 100000
rect 33782 99200 33838 100000
rect 35806 99200 35862 100000
rect 37830 99200 37886 100000
rect 39854 99200 39910 100000
rect 41878 99200 41934 100000
rect 43902 99200 43958 100000
rect 45926 99200 45982 100000
rect 47950 99200 48006 100000
rect 49974 99200 50030 100000
rect 51998 99200 52054 100000
rect 54022 99200 54078 100000
rect 56046 99200 56102 100000
rect 58070 99200 58126 100000
rect 60094 99200 60150 100000
rect 62118 99200 62174 100000
rect 64142 99200 64198 100000
rect 66166 99200 66222 100000
rect 68190 99200 68246 100000
rect 70214 99200 70270 100000
rect 72238 99200 72294 100000
rect 74262 99200 74318 100000
rect 76286 99200 76342 100000
rect 78310 99200 78366 100000
rect 80334 99200 80390 100000
rect 82358 99200 82414 100000
rect 84382 99200 84438 100000
rect 86406 99200 86462 100000
rect 88430 99200 88486 100000
rect 90454 99200 90510 100000
rect 92478 99200 92534 100000
rect 94502 99200 94558 100000
rect 96526 99200 96582 100000
rect 98550 99200 98606 100000
<< obsm2 >>
rect 1510 99144 3366 99362
rect 3534 99144 5390 99362
rect 5558 99144 7414 99362
rect 7582 99144 9438 99362
rect 9606 99144 11462 99362
rect 11630 99144 13486 99362
rect 13654 99144 15510 99362
rect 15678 99144 17534 99362
rect 17702 99144 19558 99362
rect 19726 99144 21582 99362
rect 21750 99144 23606 99362
rect 23774 99144 25630 99362
rect 25798 99144 27654 99362
rect 27822 99144 29678 99362
rect 29846 99144 31702 99362
rect 31870 99144 33726 99362
rect 33894 99144 35750 99362
rect 35918 99144 37774 99362
rect 37942 99144 39798 99362
rect 39966 99144 41822 99362
rect 41990 99144 43846 99362
rect 44014 99144 45870 99362
rect 46038 99144 47894 99362
rect 48062 99144 49918 99362
rect 50086 99144 51942 99362
rect 52110 99144 53966 99362
rect 54134 99144 55990 99362
rect 56158 99144 58014 99362
rect 58182 99144 60038 99362
rect 60206 99144 62062 99362
rect 62230 99144 64086 99362
rect 64254 99144 66110 99362
rect 66278 99144 68134 99362
rect 68302 99144 70158 99362
rect 70326 99144 72182 99362
rect 72350 99144 74206 99362
rect 74374 99144 76230 99362
rect 76398 99144 78254 99362
rect 78422 99144 80278 99362
rect 80446 99144 82302 99362
rect 82470 99144 84326 99362
rect 84494 99144 86350 99362
rect 86518 99144 88374 99362
rect 88542 99144 90398 99362
rect 90566 99144 92422 99362
rect 92590 99144 94446 99362
rect 94614 99144 96470 99362
rect 96638 99144 98494 99362
rect 1398 2139 98604 99144
<< metal3 >>
rect 99200 96568 100000 96688
rect 99200 94664 100000 94784
rect 0 92760 800 92880
rect 99200 92760 100000 92880
rect 0 91944 800 92064
rect 0 91128 800 91248
rect 99200 90856 100000 90976
rect 0 90312 800 90432
rect 0 89496 800 89616
rect 99200 88952 100000 89072
rect 0 88680 800 88800
rect 0 87864 800 87984
rect 0 87048 800 87168
rect 99200 87048 100000 87168
rect 0 86232 800 86352
rect 0 85416 800 85536
rect 99200 85144 100000 85264
rect 0 84600 800 84720
rect 0 83784 800 83904
rect 99200 83240 100000 83360
rect 0 82968 800 83088
rect 0 82152 800 82272
rect 0 81336 800 81456
rect 99200 81336 100000 81456
rect 0 80520 800 80640
rect 0 79704 800 79824
rect 99200 79432 100000 79552
rect 0 78888 800 79008
rect 0 78072 800 78192
rect 99200 77528 100000 77648
rect 0 77256 800 77376
rect 0 76440 800 76560
rect 0 75624 800 75744
rect 99200 75624 100000 75744
rect 0 74808 800 74928
rect 0 73992 800 74112
rect 99200 73720 100000 73840
rect 0 73176 800 73296
rect 0 72360 800 72480
rect 99200 71816 100000 71936
rect 0 71544 800 71664
rect 0 70728 800 70848
rect 0 69912 800 70032
rect 99200 69912 100000 70032
rect 0 69096 800 69216
rect 0 68280 800 68400
rect 99200 68008 100000 68128
rect 0 67464 800 67584
rect 0 66648 800 66768
rect 99200 66104 100000 66224
rect 0 65832 800 65952
rect 0 65016 800 65136
rect 0 64200 800 64320
rect 99200 64200 100000 64320
rect 0 63384 800 63504
rect 0 62568 800 62688
rect 99200 62296 100000 62416
rect 0 61752 800 61872
rect 0 60936 800 61056
rect 99200 60392 100000 60512
rect 0 60120 800 60240
rect 0 59304 800 59424
rect 0 58488 800 58608
rect 99200 58488 100000 58608
rect 0 57672 800 57792
rect 0 56856 800 56976
rect 99200 56584 100000 56704
rect 0 56040 800 56160
rect 0 55224 800 55344
rect 99200 54680 100000 54800
rect 0 54408 800 54528
rect 0 53592 800 53712
rect 0 52776 800 52896
rect 99200 52776 100000 52896
rect 0 51960 800 52080
rect 0 51144 800 51264
rect 99200 50872 100000 50992
rect 0 50328 800 50448
rect 0 49512 800 49632
rect 99200 48968 100000 49088
rect 0 48696 800 48816
rect 0 47880 800 48000
rect 0 47064 800 47184
rect 99200 47064 100000 47184
rect 0 46248 800 46368
rect 0 45432 800 45552
rect 99200 45160 100000 45280
rect 0 44616 800 44736
rect 0 43800 800 43920
rect 99200 43256 100000 43376
rect 0 42984 800 43104
rect 0 42168 800 42288
rect 0 41352 800 41472
rect 99200 41352 100000 41472
rect 0 40536 800 40656
rect 0 39720 800 39840
rect 99200 39448 100000 39568
rect 0 38904 800 39024
rect 0 38088 800 38208
rect 99200 37544 100000 37664
rect 0 37272 800 37392
rect 0 36456 800 36576
rect 0 35640 800 35760
rect 99200 35640 100000 35760
rect 0 34824 800 34944
rect 0 34008 800 34128
rect 99200 33736 100000 33856
rect 0 33192 800 33312
rect 0 32376 800 32496
rect 99200 31832 100000 31952
rect 0 31560 800 31680
rect 0 30744 800 30864
rect 0 29928 800 30048
rect 99200 29928 100000 30048
rect 0 29112 800 29232
rect 0 28296 800 28416
rect 99200 28024 100000 28144
rect 0 27480 800 27600
rect 0 26664 800 26784
rect 99200 26120 100000 26240
rect 0 25848 800 25968
rect 0 25032 800 25152
rect 0 24216 800 24336
rect 99200 24216 100000 24336
rect 0 23400 800 23520
rect 0 22584 800 22704
rect 99200 22312 100000 22432
rect 0 21768 800 21888
rect 0 20952 800 21072
rect 99200 20408 100000 20528
rect 0 20136 800 20256
rect 0 19320 800 19440
rect 0 18504 800 18624
rect 99200 18504 100000 18624
rect 0 17688 800 17808
rect 0 16872 800 16992
rect 99200 16600 100000 16720
rect 0 16056 800 16176
rect 0 15240 800 15360
rect 99200 14696 100000 14816
rect 0 14424 800 14544
rect 0 13608 800 13728
rect 0 12792 800 12912
rect 99200 12792 100000 12912
rect 0 11976 800 12096
rect 0 11160 800 11280
rect 99200 10888 100000 11008
rect 0 10344 800 10464
rect 0 9528 800 9648
rect 99200 8984 100000 9104
rect 0 8712 800 8832
rect 0 7896 800 8016
rect 0 7080 800 7200
rect 99200 7080 100000 7200
rect 99200 5176 100000 5296
rect 99200 3272 100000 3392
<< obsm3 >>
rect 800 96768 99200 97409
rect 800 96488 99120 96768
rect 800 94864 99200 96488
rect 800 94584 99120 94864
rect 800 92960 99200 94584
rect 880 92680 99120 92960
rect 800 92144 99200 92680
rect 880 91864 99200 92144
rect 800 91328 99200 91864
rect 880 91056 99200 91328
rect 880 91048 99120 91056
rect 800 90776 99120 91048
rect 800 90512 99200 90776
rect 880 90232 99200 90512
rect 800 89696 99200 90232
rect 880 89416 99200 89696
rect 800 89152 99200 89416
rect 800 88880 99120 89152
rect 880 88872 99120 88880
rect 880 88600 99200 88872
rect 800 88064 99200 88600
rect 880 87784 99200 88064
rect 800 87248 99200 87784
rect 880 86968 99120 87248
rect 800 86432 99200 86968
rect 880 86152 99200 86432
rect 800 85616 99200 86152
rect 880 85344 99200 85616
rect 880 85336 99120 85344
rect 800 85064 99120 85336
rect 800 84800 99200 85064
rect 880 84520 99200 84800
rect 800 83984 99200 84520
rect 880 83704 99200 83984
rect 800 83440 99200 83704
rect 800 83168 99120 83440
rect 880 83160 99120 83168
rect 880 82888 99200 83160
rect 800 82352 99200 82888
rect 880 82072 99200 82352
rect 800 81536 99200 82072
rect 880 81256 99120 81536
rect 800 80720 99200 81256
rect 880 80440 99200 80720
rect 800 79904 99200 80440
rect 880 79632 99200 79904
rect 880 79624 99120 79632
rect 800 79352 99120 79624
rect 800 79088 99200 79352
rect 880 78808 99200 79088
rect 800 78272 99200 78808
rect 880 77992 99200 78272
rect 800 77728 99200 77992
rect 800 77456 99120 77728
rect 880 77448 99120 77456
rect 880 77176 99200 77448
rect 800 76640 99200 77176
rect 880 76360 99200 76640
rect 800 75824 99200 76360
rect 880 75544 99120 75824
rect 800 75008 99200 75544
rect 880 74728 99200 75008
rect 800 74192 99200 74728
rect 880 73920 99200 74192
rect 880 73912 99120 73920
rect 800 73640 99120 73912
rect 800 73376 99200 73640
rect 880 73096 99200 73376
rect 800 72560 99200 73096
rect 880 72280 99200 72560
rect 800 72016 99200 72280
rect 800 71744 99120 72016
rect 880 71736 99120 71744
rect 880 71464 99200 71736
rect 800 70928 99200 71464
rect 880 70648 99200 70928
rect 800 70112 99200 70648
rect 880 69832 99120 70112
rect 800 69296 99200 69832
rect 880 69016 99200 69296
rect 800 68480 99200 69016
rect 880 68208 99200 68480
rect 880 68200 99120 68208
rect 800 67928 99120 68200
rect 800 67664 99200 67928
rect 880 67384 99200 67664
rect 800 66848 99200 67384
rect 880 66568 99200 66848
rect 800 66304 99200 66568
rect 800 66032 99120 66304
rect 880 66024 99120 66032
rect 880 65752 99200 66024
rect 800 65216 99200 65752
rect 880 64936 99200 65216
rect 800 64400 99200 64936
rect 880 64120 99120 64400
rect 800 63584 99200 64120
rect 880 63304 99200 63584
rect 800 62768 99200 63304
rect 880 62496 99200 62768
rect 880 62488 99120 62496
rect 800 62216 99120 62488
rect 800 61952 99200 62216
rect 880 61672 99200 61952
rect 800 61136 99200 61672
rect 880 60856 99200 61136
rect 800 60592 99200 60856
rect 800 60320 99120 60592
rect 880 60312 99120 60320
rect 880 60040 99200 60312
rect 800 59504 99200 60040
rect 880 59224 99200 59504
rect 800 58688 99200 59224
rect 880 58408 99120 58688
rect 800 57872 99200 58408
rect 880 57592 99200 57872
rect 800 57056 99200 57592
rect 880 56784 99200 57056
rect 880 56776 99120 56784
rect 800 56504 99120 56776
rect 800 56240 99200 56504
rect 880 55960 99200 56240
rect 800 55424 99200 55960
rect 880 55144 99200 55424
rect 800 54880 99200 55144
rect 800 54608 99120 54880
rect 880 54600 99120 54608
rect 880 54328 99200 54600
rect 800 53792 99200 54328
rect 880 53512 99200 53792
rect 800 52976 99200 53512
rect 880 52696 99120 52976
rect 800 52160 99200 52696
rect 880 51880 99200 52160
rect 800 51344 99200 51880
rect 880 51072 99200 51344
rect 880 51064 99120 51072
rect 800 50792 99120 51064
rect 800 50528 99200 50792
rect 880 50248 99200 50528
rect 800 49712 99200 50248
rect 880 49432 99200 49712
rect 800 49168 99200 49432
rect 800 48896 99120 49168
rect 880 48888 99120 48896
rect 880 48616 99200 48888
rect 800 48080 99200 48616
rect 880 47800 99200 48080
rect 800 47264 99200 47800
rect 880 46984 99120 47264
rect 800 46448 99200 46984
rect 880 46168 99200 46448
rect 800 45632 99200 46168
rect 880 45360 99200 45632
rect 880 45352 99120 45360
rect 800 45080 99120 45352
rect 800 44816 99200 45080
rect 880 44536 99200 44816
rect 800 44000 99200 44536
rect 880 43720 99200 44000
rect 800 43456 99200 43720
rect 800 43184 99120 43456
rect 880 43176 99120 43184
rect 880 42904 99200 43176
rect 800 42368 99200 42904
rect 880 42088 99200 42368
rect 800 41552 99200 42088
rect 880 41272 99120 41552
rect 800 40736 99200 41272
rect 880 40456 99200 40736
rect 800 39920 99200 40456
rect 880 39648 99200 39920
rect 880 39640 99120 39648
rect 800 39368 99120 39640
rect 800 39104 99200 39368
rect 880 38824 99200 39104
rect 800 38288 99200 38824
rect 880 38008 99200 38288
rect 800 37744 99200 38008
rect 800 37472 99120 37744
rect 880 37464 99120 37472
rect 880 37192 99200 37464
rect 800 36656 99200 37192
rect 880 36376 99200 36656
rect 800 35840 99200 36376
rect 880 35560 99120 35840
rect 800 35024 99200 35560
rect 880 34744 99200 35024
rect 800 34208 99200 34744
rect 880 33936 99200 34208
rect 880 33928 99120 33936
rect 800 33656 99120 33928
rect 800 33392 99200 33656
rect 880 33112 99200 33392
rect 800 32576 99200 33112
rect 880 32296 99200 32576
rect 800 32032 99200 32296
rect 800 31760 99120 32032
rect 880 31752 99120 31760
rect 880 31480 99200 31752
rect 800 30944 99200 31480
rect 880 30664 99200 30944
rect 800 30128 99200 30664
rect 880 29848 99120 30128
rect 800 29312 99200 29848
rect 880 29032 99200 29312
rect 800 28496 99200 29032
rect 880 28224 99200 28496
rect 880 28216 99120 28224
rect 800 27944 99120 28216
rect 800 27680 99200 27944
rect 880 27400 99200 27680
rect 800 26864 99200 27400
rect 880 26584 99200 26864
rect 800 26320 99200 26584
rect 800 26048 99120 26320
rect 880 26040 99120 26048
rect 880 25768 99200 26040
rect 800 25232 99200 25768
rect 880 24952 99200 25232
rect 800 24416 99200 24952
rect 880 24136 99120 24416
rect 800 23600 99200 24136
rect 880 23320 99200 23600
rect 800 22784 99200 23320
rect 880 22512 99200 22784
rect 880 22504 99120 22512
rect 800 22232 99120 22504
rect 800 21968 99200 22232
rect 880 21688 99200 21968
rect 800 21152 99200 21688
rect 880 20872 99200 21152
rect 800 20608 99200 20872
rect 800 20336 99120 20608
rect 880 20328 99120 20336
rect 880 20056 99200 20328
rect 800 19520 99200 20056
rect 880 19240 99200 19520
rect 800 18704 99200 19240
rect 880 18424 99120 18704
rect 800 17888 99200 18424
rect 880 17608 99200 17888
rect 800 17072 99200 17608
rect 880 16800 99200 17072
rect 880 16792 99120 16800
rect 800 16520 99120 16792
rect 800 16256 99200 16520
rect 880 15976 99200 16256
rect 800 15440 99200 15976
rect 880 15160 99200 15440
rect 800 14896 99200 15160
rect 800 14624 99120 14896
rect 880 14616 99120 14624
rect 880 14344 99200 14616
rect 800 13808 99200 14344
rect 880 13528 99200 13808
rect 800 12992 99200 13528
rect 880 12712 99120 12992
rect 800 12176 99200 12712
rect 880 11896 99200 12176
rect 800 11360 99200 11896
rect 880 11088 99200 11360
rect 880 11080 99120 11088
rect 800 10808 99120 11080
rect 800 10544 99200 10808
rect 880 10264 99200 10544
rect 800 9728 99200 10264
rect 880 9448 99200 9728
rect 800 9184 99200 9448
rect 800 8912 99120 9184
rect 880 8904 99120 8912
rect 880 8632 99200 8904
rect 800 8096 99200 8632
rect 880 7816 99200 8096
rect 800 7280 99200 7816
rect 880 7000 99120 7280
rect 800 5376 99200 7000
rect 800 5096 99120 5376
rect 800 3472 99200 5096
rect 800 3192 99120 3472
rect 800 2143 99200 3192
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< labels >>
rlabel metal3 s 99200 79432 100000 79552 6 addr0[0]
port 1 nsew signal output
rlabel metal3 s 99200 81336 100000 81456 6 addr0[1]
port 2 nsew signal output
rlabel metal3 s 99200 83240 100000 83360 6 addr0[2]
port 3 nsew signal output
rlabel metal3 s 99200 85144 100000 85264 6 addr0[3]
port 4 nsew signal output
rlabel metal3 s 99200 87048 100000 87168 6 addr0[4]
port 5 nsew signal output
rlabel metal3 s 99200 88952 100000 89072 6 addr0[5]
port 6 nsew signal output
rlabel metal3 s 99200 90856 100000 90976 6 addr0[6]
port 7 nsew signal output
rlabel metal3 s 99200 92760 100000 92880 6 addr0[7]
port 8 nsew signal output
rlabel metal3 s 99200 94664 100000 94784 6 addr0[8]
port 9 nsew signal output
rlabel metal3 s 99200 5176 100000 5296 6 clk0
port 10 nsew signal output
rlabel metal3 s 99200 7080 100000 7200 6 csb0
port 11 nsew signal output
rlabel metal3 s 99200 18504 100000 18624 6 din0[0]
port 12 nsew signal output
rlabel metal3 s 99200 37544 100000 37664 6 din0[10]
port 13 nsew signal output
rlabel metal3 s 99200 39448 100000 39568 6 din0[11]
port 14 nsew signal output
rlabel metal3 s 99200 41352 100000 41472 6 din0[12]
port 15 nsew signal output
rlabel metal3 s 99200 43256 100000 43376 6 din0[13]
port 16 nsew signal output
rlabel metal3 s 99200 45160 100000 45280 6 din0[14]
port 17 nsew signal output
rlabel metal3 s 99200 47064 100000 47184 6 din0[15]
port 18 nsew signal output
rlabel metal3 s 99200 48968 100000 49088 6 din0[16]
port 19 nsew signal output
rlabel metal3 s 99200 50872 100000 50992 6 din0[17]
port 20 nsew signal output
rlabel metal3 s 99200 52776 100000 52896 6 din0[18]
port 21 nsew signal output
rlabel metal3 s 99200 54680 100000 54800 6 din0[19]
port 22 nsew signal output
rlabel metal3 s 99200 20408 100000 20528 6 din0[1]
port 23 nsew signal output
rlabel metal3 s 99200 56584 100000 56704 6 din0[20]
port 24 nsew signal output
rlabel metal3 s 99200 58488 100000 58608 6 din0[21]
port 25 nsew signal output
rlabel metal3 s 99200 60392 100000 60512 6 din0[22]
port 26 nsew signal output
rlabel metal3 s 99200 62296 100000 62416 6 din0[23]
port 27 nsew signal output
rlabel metal3 s 99200 64200 100000 64320 6 din0[24]
port 28 nsew signal output
rlabel metal3 s 99200 66104 100000 66224 6 din0[25]
port 29 nsew signal output
rlabel metal3 s 99200 68008 100000 68128 6 din0[26]
port 30 nsew signal output
rlabel metal3 s 99200 69912 100000 70032 6 din0[27]
port 31 nsew signal output
rlabel metal3 s 99200 71816 100000 71936 6 din0[28]
port 32 nsew signal output
rlabel metal3 s 99200 73720 100000 73840 6 din0[29]
port 33 nsew signal output
rlabel metal3 s 99200 22312 100000 22432 6 din0[2]
port 34 nsew signal output
rlabel metal3 s 99200 75624 100000 75744 6 din0[30]
port 35 nsew signal output
rlabel metal3 s 99200 77528 100000 77648 6 din0[31]
port 36 nsew signal output
rlabel metal3 s 99200 24216 100000 24336 6 din0[3]
port 37 nsew signal output
rlabel metal3 s 99200 26120 100000 26240 6 din0[4]
port 38 nsew signal output
rlabel metal3 s 99200 28024 100000 28144 6 din0[5]
port 39 nsew signal output
rlabel metal3 s 99200 29928 100000 30048 6 din0[6]
port 40 nsew signal output
rlabel metal3 s 99200 31832 100000 31952 6 din0[7]
port 41 nsew signal output
rlabel metal3 s 99200 33736 100000 33856 6 din0[8]
port 42 nsew signal output
rlabel metal3 s 99200 35640 100000 35760 6 din0[9]
port 43 nsew signal output
rlabel metal2 s 3422 99200 3478 100000 6 dmem_addrb[0]
port 44 nsew signal input
rlabel metal2 s 9494 99200 9550 100000 6 dmem_addrb[1]
port 45 nsew signal input
rlabel metal2 s 15566 99200 15622 100000 6 dmem_addrb[2]
port 46 nsew signal input
rlabel metal2 s 21638 99200 21694 100000 6 dmem_addrb[3]
port 47 nsew signal input
rlabel metal2 s 27710 99200 27766 100000 6 dmem_addrb[4]
port 48 nsew signal input
rlabel metal2 s 33782 99200 33838 100000 6 dmem_addrb[5]
port 49 nsew signal input
rlabel metal2 s 39854 99200 39910 100000 6 dmem_addrb[6]
port 50 nsew signal input
rlabel metal2 s 45926 99200 45982 100000 6 dmem_addrb[7]
port 51 nsew signal input
rlabel metal2 s 5446 99200 5502 100000 6 dmem_addrb_o[0]
port 52 nsew signal output
rlabel metal2 s 11518 99200 11574 100000 6 dmem_addrb_o[1]
port 53 nsew signal output
rlabel metal2 s 17590 99200 17646 100000 6 dmem_addrb_o[2]
port 54 nsew signal output
rlabel metal2 s 23662 99200 23718 100000 6 dmem_addrb_o[3]
port 55 nsew signal output
rlabel metal2 s 29734 99200 29790 100000 6 dmem_addrb_o[4]
port 56 nsew signal output
rlabel metal2 s 35806 99200 35862 100000 6 dmem_addrb_o[5]
port 57 nsew signal output
rlabel metal2 s 41878 99200 41934 100000 6 dmem_addrb_o[6]
port 58 nsew signal output
rlabel metal2 s 47950 99200 48006 100000 6 dmem_addrb_o[7]
port 59 nsew signal output
rlabel metal2 s 7470 99200 7526 100000 6 dmem_doutb[0]
port 60 nsew signal input
rlabel metal2 s 56046 99200 56102 100000 6 dmem_doutb[10]
port 61 nsew signal input
rlabel metal2 s 58070 99200 58126 100000 6 dmem_doutb[11]
port 62 nsew signal input
rlabel metal2 s 60094 99200 60150 100000 6 dmem_doutb[12]
port 63 nsew signal input
rlabel metal2 s 62118 99200 62174 100000 6 dmem_doutb[13]
port 64 nsew signal input
rlabel metal2 s 64142 99200 64198 100000 6 dmem_doutb[14]
port 65 nsew signal input
rlabel metal2 s 66166 99200 66222 100000 6 dmem_doutb[15]
port 66 nsew signal input
rlabel metal2 s 68190 99200 68246 100000 6 dmem_doutb[16]
port 67 nsew signal input
rlabel metal2 s 70214 99200 70270 100000 6 dmem_doutb[17]
port 68 nsew signal input
rlabel metal2 s 72238 99200 72294 100000 6 dmem_doutb[18]
port 69 nsew signal input
rlabel metal2 s 74262 99200 74318 100000 6 dmem_doutb[19]
port 70 nsew signal input
rlabel metal2 s 13542 99200 13598 100000 6 dmem_doutb[1]
port 71 nsew signal input
rlabel metal2 s 76286 99200 76342 100000 6 dmem_doutb[20]
port 72 nsew signal input
rlabel metal2 s 78310 99200 78366 100000 6 dmem_doutb[21]
port 73 nsew signal input
rlabel metal2 s 80334 99200 80390 100000 6 dmem_doutb[22]
port 74 nsew signal input
rlabel metal2 s 82358 99200 82414 100000 6 dmem_doutb[23]
port 75 nsew signal input
rlabel metal2 s 84382 99200 84438 100000 6 dmem_doutb[24]
port 76 nsew signal input
rlabel metal2 s 86406 99200 86462 100000 6 dmem_doutb[25]
port 77 nsew signal input
rlabel metal2 s 88430 99200 88486 100000 6 dmem_doutb[26]
port 78 nsew signal input
rlabel metal2 s 90454 99200 90510 100000 6 dmem_doutb[27]
port 79 nsew signal input
rlabel metal2 s 92478 99200 92534 100000 6 dmem_doutb[28]
port 80 nsew signal input
rlabel metal2 s 94502 99200 94558 100000 6 dmem_doutb[29]
port 81 nsew signal input
rlabel metal2 s 19614 99200 19670 100000 6 dmem_doutb[2]
port 82 nsew signal input
rlabel metal2 s 96526 99200 96582 100000 6 dmem_doutb[30]
port 83 nsew signal input
rlabel metal2 s 98550 99200 98606 100000 6 dmem_doutb[31]
port 84 nsew signal input
rlabel metal2 s 25686 99200 25742 100000 6 dmem_doutb[3]
port 85 nsew signal input
rlabel metal2 s 31758 99200 31814 100000 6 dmem_doutb[4]
port 86 nsew signal input
rlabel metal2 s 37830 99200 37886 100000 6 dmem_doutb[5]
port 87 nsew signal input
rlabel metal2 s 43902 99200 43958 100000 6 dmem_doutb[6]
port 88 nsew signal input
rlabel metal2 s 49974 99200 50030 100000 6 dmem_doutb[7]
port 89 nsew signal input
rlabel metal2 s 51998 99200 52054 100000 6 dmem_doutb[8]
port 90 nsew signal input
rlabel metal2 s 54022 99200 54078 100000 6 dmem_doutb[9]
port 91 nsew signal input
rlabel metal2 s 1398 99200 1454 100000 6 dmem_enb
port 92 nsew signal input
rlabel metal3 s 99200 3272 100000 3392 6 imem_rd_cs1
port 93 nsew signal output
rlabel metal3 s 99200 96568 100000 96688 6 processor_reset
port 94 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 95 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 95 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 95 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 95 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 96 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 96 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 96 nsew ground bidirectional
rlabel metal3 s 0 7080 800 7200 6 wb_clk_i
port 97 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 wb_rst_i
port 98 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 wbs_ack_o
port 99 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 wbs_adr_i[0]
port 100 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 wbs_adr_i[10]
port 101 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 wbs_adr_i[11]
port 102 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 wbs_adr_i[12]
port 103 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 wbs_adr_i[13]
port 104 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 wbs_adr_i[14]
port 105 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 wbs_adr_i[15]
port 106 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 wbs_adr_i[16]
port 107 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 wbs_adr_i[17]
port 108 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 wbs_adr_i[18]
port 109 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 wbs_adr_i[19]
port 110 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 wbs_adr_i[1]
port 111 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 wbs_adr_i[20]
port 112 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 wbs_adr_i[21]
port 113 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 wbs_adr_i[22]
port 114 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 wbs_adr_i[23]
port 115 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 wbs_adr_i[24]
port 116 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 wbs_adr_i[25]
port 117 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 wbs_adr_i[26]
port 118 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 wbs_adr_i[27]
port 119 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 wbs_adr_i[28]
port 120 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 wbs_adr_i[29]
port 121 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 wbs_adr_i[2]
port 122 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 wbs_adr_i[30]
port 123 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 wbs_adr_i[31]
port 124 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 wbs_adr_i[3]
port 125 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 wbs_adr_i[4]
port 126 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wbs_adr_i[5]
port 127 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 wbs_adr_i[6]
port 128 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 wbs_adr_i[7]
port 129 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 wbs_adr_i[8]
port 130 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 wbs_adr_i[9]
port 131 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wbs_cyc_i
port 132 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 wbs_dat_i[0]
port 133 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 wbs_dat_i[10]
port 134 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 wbs_dat_i[11]
port 135 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 wbs_dat_i[12]
port 136 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 wbs_dat_i[13]
port 137 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 wbs_dat_i[14]
port 138 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 wbs_dat_i[15]
port 139 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 wbs_dat_i[16]
port 140 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 wbs_dat_i[17]
port 141 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 wbs_dat_i[18]
port 142 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 wbs_dat_i[19]
port 143 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 wbs_dat_i[1]
port 144 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 wbs_dat_i[20]
port 145 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 wbs_dat_i[21]
port 146 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 wbs_dat_i[22]
port 147 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbs_dat_i[23]
port 148 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 wbs_dat_i[24]
port 149 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 wbs_dat_i[25]
port 150 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 wbs_dat_i[26]
port 151 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 wbs_dat_i[27]
port 152 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 wbs_dat_i[28]
port 153 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 wbs_dat_i[29]
port 154 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 wbs_dat_i[2]
port 155 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 wbs_dat_i[30]
port 156 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 wbs_dat_i[31]
port 157 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 wbs_dat_i[3]
port 158 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_dat_i[4]
port 159 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 wbs_dat_i[5]
port 160 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wbs_dat_i[6]
port 161 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 wbs_dat_i[7]
port 162 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 wbs_dat_i[8]
port 163 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 wbs_dat_i[9]
port 164 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 wbs_dat_o[0]
port 165 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 wbs_dat_o[10]
port 166 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 wbs_dat_o[11]
port 167 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 wbs_dat_o[12]
port 168 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 wbs_dat_o[13]
port 169 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 wbs_dat_o[14]
port 170 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 wbs_dat_o[15]
port 171 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 wbs_dat_o[16]
port 172 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 wbs_dat_o[17]
port 173 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 wbs_dat_o[18]
port 174 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 wbs_dat_o[19]
port 175 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 wbs_dat_o[1]
port 176 nsew signal output
rlabel metal3 s 0 65832 800 65952 6 wbs_dat_o[20]
port 177 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 wbs_dat_o[21]
port 178 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 wbs_dat_o[22]
port 179 nsew signal output
rlabel metal3 s 0 73176 800 73296 6 wbs_dat_o[23]
port 180 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 wbs_dat_o[24]
port 181 nsew signal output
rlabel metal3 s 0 78072 800 78192 6 wbs_dat_o[25]
port 182 nsew signal output
rlabel metal3 s 0 80520 800 80640 6 wbs_dat_o[26]
port 183 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 wbs_dat_o[27]
port 184 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 wbs_dat_o[28]
port 185 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 wbs_dat_o[29]
port 186 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 wbs_dat_o[2]
port 187 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 wbs_dat_o[30]
port 188 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 wbs_dat_o[31]
port 189 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 wbs_dat_o[3]
port 190 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 wbs_dat_o[4]
port 191 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 wbs_dat_o[5]
port 192 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 wbs_dat_o[6]
port 193 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 wbs_dat_o[7]
port 194 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 wbs_dat_o[8]
port 195 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 wbs_dat_o[9]
port 196 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 wbs_sel_i[0]
port 197 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wbs_sel_i[1]
port 198 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 wbs_sel_i[2]
port 199 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 wbs_sel_i[3]
port 200 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 wbs_stb_i
port 201 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 wbs_we_i
port 202 nsew signal input
rlabel metal3 s 99200 8984 100000 9104 6 web0
port 203 nsew signal output
rlabel metal3 s 99200 10888 100000 11008 6 wmask0[0]
port 204 nsew signal output
rlabel metal3 s 99200 12792 100000 12912 6 wmask0[1]
port 205 nsew signal output
rlabel metal3 s 99200 14696 100000 14816 6 wmask0[2]
port 206 nsew signal output
rlabel metal3 s 99200 16600 100000 16720 6 wmask0[3]
port 207 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3281562
string GDS_FILE /home/ali11-2000/efabless/mpw-waprv/openlane/wb_interface/runs/22_09_11_17_12/results/signoff/wb_interface.magic.gds
string GDS_START 150022
<< end >>

