magic
tech sky130B
magscale 1 2
timestamp 1662897243
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 484 178848 118924
<< metal2 >>
rect 3054 119200 3110 120000
rect 5814 119200 5870 120000
rect 8574 119200 8630 120000
rect 11334 119200 11390 120000
rect 14094 119200 14150 120000
rect 16854 119200 16910 120000
rect 19614 119200 19670 120000
rect 22374 119200 22430 120000
rect 25134 119200 25190 120000
rect 27894 119200 27950 120000
rect 30654 119200 30710 120000
rect 33414 119200 33470 120000
rect 36174 119200 36230 120000
rect 38934 119200 38990 120000
rect 41694 119200 41750 120000
rect 44454 119200 44510 120000
rect 47214 119200 47270 120000
rect 49974 119200 50030 120000
rect 52734 119200 52790 120000
rect 55494 119200 55550 120000
rect 58254 119200 58310 120000
rect 61014 119200 61070 120000
rect 63774 119200 63830 120000
rect 66534 119200 66590 120000
rect 69294 119200 69350 120000
rect 72054 119200 72110 120000
rect 74814 119200 74870 120000
rect 77574 119200 77630 120000
rect 80334 119200 80390 120000
rect 83094 119200 83150 120000
rect 85854 119200 85910 120000
rect 88614 119200 88670 120000
rect 91374 119200 91430 120000
rect 94134 119200 94190 120000
rect 96894 119200 96950 120000
rect 99654 119200 99710 120000
rect 102414 119200 102470 120000
rect 105174 119200 105230 120000
rect 107934 119200 107990 120000
rect 110694 119200 110750 120000
rect 113454 119200 113510 120000
rect 116214 119200 116270 120000
rect 118974 119200 119030 120000
rect 121734 119200 121790 120000
rect 124494 119200 124550 120000
rect 127254 119200 127310 120000
rect 130014 119200 130070 120000
rect 132774 119200 132830 120000
rect 135534 119200 135590 120000
rect 138294 119200 138350 120000
rect 141054 119200 141110 120000
rect 143814 119200 143870 120000
rect 146574 119200 146630 120000
rect 149334 119200 149390 120000
rect 152094 119200 152150 120000
rect 154854 119200 154910 120000
rect 157614 119200 157670 120000
rect 160374 119200 160430 120000
rect 163134 119200 163190 120000
rect 165894 119200 165950 120000
rect 168654 119200 168710 120000
rect 171414 119200 171470 120000
rect 174174 119200 174230 120000
rect 176934 119200 176990 120000
rect 3054 0 3110 800
rect 5814 0 5870 800
rect 8574 0 8630 800
rect 11334 0 11390 800
rect 14094 0 14150 800
rect 16854 0 16910 800
rect 19614 0 19670 800
rect 22374 0 22430 800
rect 25134 0 25190 800
rect 27894 0 27950 800
rect 30654 0 30710 800
rect 33414 0 33470 800
rect 36174 0 36230 800
rect 38934 0 38990 800
rect 41694 0 41750 800
rect 44454 0 44510 800
rect 47214 0 47270 800
rect 49974 0 50030 800
rect 52734 0 52790 800
rect 55494 0 55550 800
rect 58254 0 58310 800
rect 61014 0 61070 800
rect 63774 0 63830 800
rect 66534 0 66590 800
rect 69294 0 69350 800
rect 72054 0 72110 800
rect 74814 0 74870 800
rect 77574 0 77630 800
rect 80334 0 80390 800
rect 83094 0 83150 800
rect 85854 0 85910 800
rect 88614 0 88670 800
rect 91374 0 91430 800
rect 94134 0 94190 800
rect 96894 0 96950 800
rect 99654 0 99710 800
rect 102414 0 102470 800
rect 105174 0 105230 800
rect 107934 0 107990 800
rect 110694 0 110750 800
rect 113454 0 113510 800
rect 116214 0 116270 800
rect 118974 0 119030 800
rect 121734 0 121790 800
rect 124494 0 124550 800
rect 127254 0 127310 800
rect 130014 0 130070 800
rect 132774 0 132830 800
rect 135534 0 135590 800
rect 138294 0 138350 800
rect 141054 0 141110 800
rect 143814 0 143870 800
rect 146574 0 146630 800
rect 149334 0 149390 800
rect 152094 0 152150 800
rect 154854 0 154910 800
rect 157614 0 157670 800
rect 160374 0 160430 800
rect 163134 0 163190 800
rect 165894 0 165950 800
rect 168654 0 168710 800
rect 171414 0 171470 800
rect 174174 0 174230 800
rect 176934 0 176990 800
<< obsm2 >>
rect 1398 119144 2998 119354
rect 3166 119144 5758 119354
rect 5926 119144 8518 119354
rect 8686 119144 11278 119354
rect 11446 119144 14038 119354
rect 14206 119144 16798 119354
rect 16966 119144 19558 119354
rect 19726 119144 22318 119354
rect 22486 119144 25078 119354
rect 25246 119144 27838 119354
rect 28006 119144 30598 119354
rect 30766 119144 33358 119354
rect 33526 119144 36118 119354
rect 36286 119144 38878 119354
rect 39046 119144 41638 119354
rect 41806 119144 44398 119354
rect 44566 119144 47158 119354
rect 47326 119144 49918 119354
rect 50086 119144 52678 119354
rect 52846 119144 55438 119354
rect 55606 119144 58198 119354
rect 58366 119144 60958 119354
rect 61126 119144 63718 119354
rect 63886 119144 66478 119354
rect 66646 119144 69238 119354
rect 69406 119144 71998 119354
rect 72166 119144 74758 119354
rect 74926 119144 77518 119354
rect 77686 119144 80278 119354
rect 80446 119144 83038 119354
rect 83206 119144 85798 119354
rect 85966 119144 88558 119354
rect 88726 119144 91318 119354
rect 91486 119144 94078 119354
rect 94246 119144 96838 119354
rect 97006 119144 99598 119354
rect 99766 119144 102358 119354
rect 102526 119144 105118 119354
rect 105286 119144 107878 119354
rect 108046 119144 110638 119354
rect 110806 119144 113398 119354
rect 113566 119144 116158 119354
rect 116326 119144 118918 119354
rect 119086 119144 121678 119354
rect 121846 119144 124438 119354
rect 124606 119144 127198 119354
rect 127366 119144 129958 119354
rect 130126 119144 132718 119354
rect 132886 119144 135478 119354
rect 135646 119144 138238 119354
rect 138406 119144 140998 119354
rect 141166 119144 143758 119354
rect 143926 119144 146518 119354
rect 146686 119144 149278 119354
rect 149446 119144 152038 119354
rect 152206 119144 154798 119354
rect 154966 119144 157558 119354
rect 157726 119144 160318 119354
rect 160486 119144 163078 119354
rect 163246 119144 165838 119354
rect 166006 119144 168598 119354
rect 168766 119144 171358 119354
rect 171526 119144 174118 119354
rect 174286 119144 176878 119354
rect 177046 119144 178644 119354
rect 1398 856 178644 119144
rect 1398 478 2998 856
rect 3166 478 5758 856
rect 5926 478 8518 856
rect 8686 478 11278 856
rect 11446 478 14038 856
rect 14206 478 16798 856
rect 16966 478 19558 856
rect 19726 478 22318 856
rect 22486 478 25078 856
rect 25246 478 27838 856
rect 28006 478 30598 856
rect 30766 478 33358 856
rect 33526 478 36118 856
rect 36286 478 38878 856
rect 39046 478 41638 856
rect 41806 478 44398 856
rect 44566 478 47158 856
rect 47326 478 49918 856
rect 50086 478 52678 856
rect 52846 478 55438 856
rect 55606 478 58198 856
rect 58366 478 60958 856
rect 61126 478 63718 856
rect 63886 478 66478 856
rect 66646 478 69238 856
rect 69406 478 71998 856
rect 72166 478 74758 856
rect 74926 478 77518 856
rect 77686 478 80278 856
rect 80446 478 83038 856
rect 83206 478 85798 856
rect 85966 478 88558 856
rect 88726 478 91318 856
rect 91486 478 94078 856
rect 94246 478 96838 856
rect 97006 478 99598 856
rect 99766 478 102358 856
rect 102526 478 105118 856
rect 105286 478 107878 856
rect 108046 478 110638 856
rect 110806 478 113398 856
rect 113566 478 116158 856
rect 116326 478 118918 856
rect 119086 478 121678 856
rect 121846 478 124438 856
rect 124606 478 127198 856
rect 127366 478 129958 856
rect 130126 478 132718 856
rect 132886 478 135478 856
rect 135646 478 138238 856
rect 138406 478 140998 856
rect 141166 478 143758 856
rect 143926 478 146518 856
rect 146686 478 149278 856
rect 149446 478 152038 856
rect 152206 478 154798 856
rect 154966 478 157558 856
rect 157726 478 160318 856
rect 160486 478 163078 856
rect 163246 478 165838 856
rect 166006 478 168598 856
rect 168766 478 171358 856
rect 171526 478 174118 856
rect 174286 478 176878 856
rect 177046 478 178644 856
<< metal3 >>
rect 0 116016 800 116136
rect 179200 115200 180000 115320
rect 179200 113704 180000 113824
rect 0 112616 800 112736
rect 179200 112208 180000 112328
rect 179200 110712 180000 110832
rect 0 109216 800 109336
rect 179200 109216 180000 109336
rect 179200 107720 180000 107840
rect 179200 106224 180000 106344
rect 0 105816 800 105936
rect 179200 104728 180000 104848
rect 179200 103232 180000 103352
rect 0 102416 800 102536
rect 179200 101736 180000 101856
rect 179200 100240 180000 100360
rect 0 99016 800 99136
rect 179200 98744 180000 98864
rect 179200 97248 180000 97368
rect 0 95616 800 95736
rect 179200 95752 180000 95872
rect 179200 94256 180000 94376
rect 179200 92760 180000 92880
rect 0 92216 800 92336
rect 179200 91264 180000 91384
rect 179200 89768 180000 89888
rect 0 88816 800 88936
rect 179200 88272 180000 88392
rect 179200 86776 180000 86896
rect 0 85416 800 85536
rect 179200 85280 180000 85400
rect 179200 83784 180000 83904
rect 179200 82288 180000 82408
rect 0 82016 800 82136
rect 179200 80792 180000 80912
rect 179200 79296 180000 79416
rect 0 78616 800 78736
rect 179200 77800 180000 77920
rect 179200 76304 180000 76424
rect 0 75216 800 75336
rect 179200 74808 180000 74928
rect 179200 73312 180000 73432
rect 0 71816 800 71936
rect 179200 71816 180000 71936
rect 179200 70320 180000 70440
rect 179200 68824 180000 68944
rect 0 68416 800 68536
rect 179200 67328 180000 67448
rect 179200 65832 180000 65952
rect 0 65016 800 65136
rect 179200 64336 180000 64456
rect 179200 62840 180000 62960
rect 0 61616 800 61736
rect 179200 61344 180000 61464
rect 179200 59848 180000 59968
rect 0 58216 800 58336
rect 179200 58352 180000 58472
rect 179200 56856 180000 56976
rect 179200 55360 180000 55480
rect 0 54816 800 54936
rect 179200 53864 180000 53984
rect 179200 52368 180000 52488
rect 0 51416 800 51536
rect 179200 50872 180000 50992
rect 179200 49376 180000 49496
rect 0 48016 800 48136
rect 179200 47880 180000 48000
rect 179200 46384 180000 46504
rect 179200 44888 180000 45008
rect 0 44616 800 44736
rect 179200 43392 180000 43512
rect 179200 41896 180000 42016
rect 0 41216 800 41336
rect 179200 40400 180000 40520
rect 179200 38904 180000 39024
rect 0 37816 800 37936
rect 179200 37408 180000 37528
rect 179200 35912 180000 36032
rect 0 34416 800 34536
rect 179200 34416 180000 34536
rect 179200 32920 180000 33040
rect 179200 31424 180000 31544
rect 0 31016 800 31136
rect 179200 29928 180000 30048
rect 179200 28432 180000 28552
rect 0 27616 800 27736
rect 179200 26936 180000 27056
rect 179200 25440 180000 25560
rect 0 24216 800 24336
rect 179200 23944 180000 24064
rect 179200 22448 180000 22568
rect 0 20816 800 20936
rect 179200 20952 180000 21072
rect 179200 19456 180000 19576
rect 179200 17960 180000 18080
rect 0 17416 800 17536
rect 179200 16464 180000 16584
rect 179200 14968 180000 15088
rect 0 14016 800 14136
rect 179200 13472 180000 13592
rect 179200 11976 180000 12096
rect 0 10616 800 10736
rect 179200 10480 180000 10600
rect 179200 8984 180000 9104
rect 179200 7488 180000 7608
rect 0 7216 800 7336
rect 179200 5992 180000 6112
rect 179200 4496 180000 4616
rect 0 3816 800 3936
<< obsm3 >>
rect 800 116216 179200 117537
rect 880 115936 179200 116216
rect 800 115400 179200 115936
rect 800 115120 179120 115400
rect 800 113904 179200 115120
rect 800 113624 179120 113904
rect 800 112816 179200 113624
rect 880 112536 179200 112816
rect 800 112408 179200 112536
rect 800 112128 179120 112408
rect 800 110912 179200 112128
rect 800 110632 179120 110912
rect 800 109416 179200 110632
rect 880 109136 179120 109416
rect 800 107920 179200 109136
rect 800 107640 179120 107920
rect 800 106424 179200 107640
rect 800 106144 179120 106424
rect 800 106016 179200 106144
rect 880 105736 179200 106016
rect 800 104928 179200 105736
rect 800 104648 179120 104928
rect 800 103432 179200 104648
rect 800 103152 179120 103432
rect 800 102616 179200 103152
rect 880 102336 179200 102616
rect 800 101936 179200 102336
rect 800 101656 179120 101936
rect 800 100440 179200 101656
rect 800 100160 179120 100440
rect 800 99216 179200 100160
rect 880 98944 179200 99216
rect 880 98936 179120 98944
rect 800 98664 179120 98936
rect 800 97448 179200 98664
rect 800 97168 179120 97448
rect 800 95952 179200 97168
rect 800 95816 179120 95952
rect 880 95672 179120 95816
rect 880 95536 179200 95672
rect 800 94456 179200 95536
rect 800 94176 179120 94456
rect 800 92960 179200 94176
rect 800 92680 179120 92960
rect 800 92416 179200 92680
rect 880 92136 179200 92416
rect 800 91464 179200 92136
rect 800 91184 179120 91464
rect 800 89968 179200 91184
rect 800 89688 179120 89968
rect 800 89016 179200 89688
rect 880 88736 179200 89016
rect 800 88472 179200 88736
rect 800 88192 179120 88472
rect 800 86976 179200 88192
rect 800 86696 179120 86976
rect 800 85616 179200 86696
rect 880 85480 179200 85616
rect 880 85336 179120 85480
rect 800 85200 179120 85336
rect 800 83984 179200 85200
rect 800 83704 179120 83984
rect 800 82488 179200 83704
rect 800 82216 179120 82488
rect 880 82208 179120 82216
rect 880 81936 179200 82208
rect 800 80992 179200 81936
rect 800 80712 179120 80992
rect 800 79496 179200 80712
rect 800 79216 179120 79496
rect 800 78816 179200 79216
rect 880 78536 179200 78816
rect 800 78000 179200 78536
rect 800 77720 179120 78000
rect 800 76504 179200 77720
rect 800 76224 179120 76504
rect 800 75416 179200 76224
rect 880 75136 179200 75416
rect 800 75008 179200 75136
rect 800 74728 179120 75008
rect 800 73512 179200 74728
rect 800 73232 179120 73512
rect 800 72016 179200 73232
rect 880 71736 179120 72016
rect 800 70520 179200 71736
rect 800 70240 179120 70520
rect 800 69024 179200 70240
rect 800 68744 179120 69024
rect 800 68616 179200 68744
rect 880 68336 179200 68616
rect 800 67528 179200 68336
rect 800 67248 179120 67528
rect 800 66032 179200 67248
rect 800 65752 179120 66032
rect 800 65216 179200 65752
rect 880 64936 179200 65216
rect 800 64536 179200 64936
rect 800 64256 179120 64536
rect 800 63040 179200 64256
rect 800 62760 179120 63040
rect 800 61816 179200 62760
rect 880 61544 179200 61816
rect 880 61536 179120 61544
rect 800 61264 179120 61536
rect 800 60048 179200 61264
rect 800 59768 179120 60048
rect 800 58552 179200 59768
rect 800 58416 179120 58552
rect 880 58272 179120 58416
rect 880 58136 179200 58272
rect 800 57056 179200 58136
rect 800 56776 179120 57056
rect 800 55560 179200 56776
rect 800 55280 179120 55560
rect 800 55016 179200 55280
rect 880 54736 179200 55016
rect 800 54064 179200 54736
rect 800 53784 179120 54064
rect 800 52568 179200 53784
rect 800 52288 179120 52568
rect 800 51616 179200 52288
rect 880 51336 179200 51616
rect 800 51072 179200 51336
rect 800 50792 179120 51072
rect 800 49576 179200 50792
rect 800 49296 179120 49576
rect 800 48216 179200 49296
rect 880 48080 179200 48216
rect 880 47936 179120 48080
rect 800 47800 179120 47936
rect 800 46584 179200 47800
rect 800 46304 179120 46584
rect 800 45088 179200 46304
rect 800 44816 179120 45088
rect 880 44808 179120 44816
rect 880 44536 179200 44808
rect 800 43592 179200 44536
rect 800 43312 179120 43592
rect 800 42096 179200 43312
rect 800 41816 179120 42096
rect 800 41416 179200 41816
rect 880 41136 179200 41416
rect 800 40600 179200 41136
rect 800 40320 179120 40600
rect 800 39104 179200 40320
rect 800 38824 179120 39104
rect 800 38016 179200 38824
rect 880 37736 179200 38016
rect 800 37608 179200 37736
rect 800 37328 179120 37608
rect 800 36112 179200 37328
rect 800 35832 179120 36112
rect 800 34616 179200 35832
rect 880 34336 179120 34616
rect 800 33120 179200 34336
rect 800 32840 179120 33120
rect 800 31624 179200 32840
rect 800 31344 179120 31624
rect 800 31216 179200 31344
rect 880 30936 179200 31216
rect 800 30128 179200 30936
rect 800 29848 179120 30128
rect 800 28632 179200 29848
rect 800 28352 179120 28632
rect 800 27816 179200 28352
rect 880 27536 179200 27816
rect 800 27136 179200 27536
rect 800 26856 179120 27136
rect 800 25640 179200 26856
rect 800 25360 179120 25640
rect 800 24416 179200 25360
rect 880 24144 179200 24416
rect 880 24136 179120 24144
rect 800 23864 179120 24136
rect 800 22648 179200 23864
rect 800 22368 179120 22648
rect 800 21152 179200 22368
rect 800 21016 179120 21152
rect 880 20872 179120 21016
rect 880 20736 179200 20872
rect 800 19656 179200 20736
rect 800 19376 179120 19656
rect 800 18160 179200 19376
rect 800 17880 179120 18160
rect 800 17616 179200 17880
rect 880 17336 179200 17616
rect 800 16664 179200 17336
rect 800 16384 179120 16664
rect 800 15168 179200 16384
rect 800 14888 179120 15168
rect 800 14216 179200 14888
rect 880 13936 179200 14216
rect 800 13672 179200 13936
rect 800 13392 179120 13672
rect 800 12176 179200 13392
rect 800 11896 179120 12176
rect 800 10816 179200 11896
rect 880 10680 179200 10816
rect 880 10536 179120 10680
rect 800 10400 179120 10536
rect 800 9184 179200 10400
rect 800 8904 179120 9184
rect 800 7688 179200 8904
rect 800 7416 179120 7688
rect 880 7408 179120 7416
rect 880 7136 179200 7408
rect 800 6192 179200 7136
rect 800 5912 179120 6192
rect 800 4696 179200 5912
rect 800 4416 179120 4696
rect 800 4016 179200 4416
rect 880 3736 179200 4016
rect 800 716 179200 3736
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 9443 2048 19488 116517
rect 19968 2048 34848 116517
rect 35328 2048 50208 116517
rect 50688 2048 65568 116517
rect 66048 2048 80928 116517
rect 81408 2048 96288 116517
rect 96768 2048 111648 116517
rect 112128 2048 127008 116517
rect 127488 2048 142368 116517
rect 142848 2048 157728 116517
rect 158208 2048 173088 116517
rect 173568 2048 177869 116517
rect 9443 715 177869 2048
<< labels >>
rlabel metal3 s 0 3816 800 3936 6 clk
port 1 nsew signal input
rlabel metal2 s 3054 119200 3110 120000 6 dmem_addra[0]
port 2 nsew signal output
rlabel metal2 s 30654 119200 30710 120000 6 dmem_addra[10]
port 3 nsew signal output
rlabel metal2 s 33414 119200 33470 120000 6 dmem_addra[11]
port 4 nsew signal output
rlabel metal2 s 36174 119200 36230 120000 6 dmem_addra[12]
port 5 nsew signal output
rlabel metal2 s 38934 119200 38990 120000 6 dmem_addra[13]
port 6 nsew signal output
rlabel metal2 s 41694 119200 41750 120000 6 dmem_addra[14]
port 7 nsew signal output
rlabel metal2 s 44454 119200 44510 120000 6 dmem_addra[15]
port 8 nsew signal output
rlabel metal2 s 47214 119200 47270 120000 6 dmem_addra[16]
port 9 nsew signal output
rlabel metal2 s 49974 119200 50030 120000 6 dmem_addra[17]
port 10 nsew signal output
rlabel metal2 s 52734 119200 52790 120000 6 dmem_addra[18]
port 11 nsew signal output
rlabel metal2 s 55494 119200 55550 120000 6 dmem_addra[19]
port 12 nsew signal output
rlabel metal2 s 5814 119200 5870 120000 6 dmem_addra[1]
port 13 nsew signal output
rlabel metal2 s 58254 119200 58310 120000 6 dmem_addra[20]
port 14 nsew signal output
rlabel metal2 s 61014 119200 61070 120000 6 dmem_addra[21]
port 15 nsew signal output
rlabel metal2 s 63774 119200 63830 120000 6 dmem_addra[22]
port 16 nsew signal output
rlabel metal2 s 66534 119200 66590 120000 6 dmem_addra[23]
port 17 nsew signal output
rlabel metal2 s 69294 119200 69350 120000 6 dmem_addra[24]
port 18 nsew signal output
rlabel metal2 s 72054 119200 72110 120000 6 dmem_addra[25]
port 19 nsew signal output
rlabel metal2 s 74814 119200 74870 120000 6 dmem_addra[26]
port 20 nsew signal output
rlabel metal2 s 77574 119200 77630 120000 6 dmem_addra[27]
port 21 nsew signal output
rlabel metal2 s 80334 119200 80390 120000 6 dmem_addra[28]
port 22 nsew signal output
rlabel metal2 s 83094 119200 83150 120000 6 dmem_addra[29]
port 23 nsew signal output
rlabel metal2 s 8574 119200 8630 120000 6 dmem_addra[2]
port 24 nsew signal output
rlabel metal2 s 85854 119200 85910 120000 6 dmem_addra[30]
port 25 nsew signal output
rlabel metal2 s 88614 119200 88670 120000 6 dmem_addra[31]
port 26 nsew signal output
rlabel metal2 s 11334 119200 11390 120000 6 dmem_addra[3]
port 27 nsew signal output
rlabel metal2 s 14094 119200 14150 120000 6 dmem_addra[4]
port 28 nsew signal output
rlabel metal2 s 16854 119200 16910 120000 6 dmem_addra[5]
port 29 nsew signal output
rlabel metal2 s 19614 119200 19670 120000 6 dmem_addra[6]
port 30 nsew signal output
rlabel metal2 s 22374 119200 22430 120000 6 dmem_addra[7]
port 31 nsew signal output
rlabel metal2 s 25134 119200 25190 120000 6 dmem_addra[8]
port 32 nsew signal output
rlabel metal2 s 27894 119200 27950 120000 6 dmem_addra[9]
port 33 nsew signal output
rlabel metal2 s 91374 119200 91430 120000 6 dmem_addrb[0]
port 34 nsew signal output
rlabel metal2 s 118974 119200 119030 120000 6 dmem_addrb[10]
port 35 nsew signal output
rlabel metal2 s 121734 119200 121790 120000 6 dmem_addrb[11]
port 36 nsew signal output
rlabel metal2 s 124494 119200 124550 120000 6 dmem_addrb[12]
port 37 nsew signal output
rlabel metal2 s 127254 119200 127310 120000 6 dmem_addrb[13]
port 38 nsew signal output
rlabel metal2 s 130014 119200 130070 120000 6 dmem_addrb[14]
port 39 nsew signal output
rlabel metal2 s 132774 119200 132830 120000 6 dmem_addrb[15]
port 40 nsew signal output
rlabel metal2 s 135534 119200 135590 120000 6 dmem_addrb[16]
port 41 nsew signal output
rlabel metal2 s 138294 119200 138350 120000 6 dmem_addrb[17]
port 42 nsew signal output
rlabel metal2 s 141054 119200 141110 120000 6 dmem_addrb[18]
port 43 nsew signal output
rlabel metal2 s 143814 119200 143870 120000 6 dmem_addrb[19]
port 44 nsew signal output
rlabel metal2 s 94134 119200 94190 120000 6 dmem_addrb[1]
port 45 nsew signal output
rlabel metal2 s 146574 119200 146630 120000 6 dmem_addrb[20]
port 46 nsew signal output
rlabel metal2 s 149334 119200 149390 120000 6 dmem_addrb[21]
port 47 nsew signal output
rlabel metal2 s 152094 119200 152150 120000 6 dmem_addrb[22]
port 48 nsew signal output
rlabel metal2 s 154854 119200 154910 120000 6 dmem_addrb[23]
port 49 nsew signal output
rlabel metal2 s 157614 119200 157670 120000 6 dmem_addrb[24]
port 50 nsew signal output
rlabel metal2 s 160374 119200 160430 120000 6 dmem_addrb[25]
port 51 nsew signal output
rlabel metal2 s 163134 119200 163190 120000 6 dmem_addrb[26]
port 52 nsew signal output
rlabel metal2 s 165894 119200 165950 120000 6 dmem_addrb[27]
port 53 nsew signal output
rlabel metal2 s 168654 119200 168710 120000 6 dmem_addrb[28]
port 54 nsew signal output
rlabel metal2 s 171414 119200 171470 120000 6 dmem_addrb[29]
port 55 nsew signal output
rlabel metal2 s 96894 119200 96950 120000 6 dmem_addrb[2]
port 56 nsew signal output
rlabel metal2 s 174174 119200 174230 120000 6 dmem_addrb[30]
port 57 nsew signal output
rlabel metal2 s 176934 119200 176990 120000 6 dmem_addrb[31]
port 58 nsew signal output
rlabel metal2 s 99654 119200 99710 120000 6 dmem_addrb[3]
port 59 nsew signal output
rlabel metal2 s 102414 119200 102470 120000 6 dmem_addrb[4]
port 60 nsew signal output
rlabel metal2 s 105174 119200 105230 120000 6 dmem_addrb[5]
port 61 nsew signal output
rlabel metal2 s 107934 119200 107990 120000 6 dmem_addrb[6]
port 62 nsew signal output
rlabel metal2 s 110694 119200 110750 120000 6 dmem_addrb[7]
port 63 nsew signal output
rlabel metal2 s 113454 119200 113510 120000 6 dmem_addrb[8]
port 64 nsew signal output
rlabel metal2 s 116214 119200 116270 120000 6 dmem_addrb[9]
port 65 nsew signal output
rlabel metal3 s 179200 4496 180000 4616 6 dmem_dina[0]
port 66 nsew signal output
rlabel metal3 s 179200 19456 180000 19576 6 dmem_dina[10]
port 67 nsew signal output
rlabel metal3 s 179200 20952 180000 21072 6 dmem_dina[11]
port 68 nsew signal output
rlabel metal3 s 179200 22448 180000 22568 6 dmem_dina[12]
port 69 nsew signal output
rlabel metal3 s 179200 23944 180000 24064 6 dmem_dina[13]
port 70 nsew signal output
rlabel metal3 s 179200 25440 180000 25560 6 dmem_dina[14]
port 71 nsew signal output
rlabel metal3 s 179200 26936 180000 27056 6 dmem_dina[15]
port 72 nsew signal output
rlabel metal3 s 179200 28432 180000 28552 6 dmem_dina[16]
port 73 nsew signal output
rlabel metal3 s 179200 29928 180000 30048 6 dmem_dina[17]
port 74 nsew signal output
rlabel metal3 s 179200 31424 180000 31544 6 dmem_dina[18]
port 75 nsew signal output
rlabel metal3 s 179200 32920 180000 33040 6 dmem_dina[19]
port 76 nsew signal output
rlabel metal3 s 179200 5992 180000 6112 6 dmem_dina[1]
port 77 nsew signal output
rlabel metal3 s 179200 34416 180000 34536 6 dmem_dina[20]
port 78 nsew signal output
rlabel metal3 s 179200 35912 180000 36032 6 dmem_dina[21]
port 79 nsew signal output
rlabel metal3 s 179200 37408 180000 37528 6 dmem_dina[22]
port 80 nsew signal output
rlabel metal3 s 179200 38904 180000 39024 6 dmem_dina[23]
port 81 nsew signal output
rlabel metal3 s 179200 40400 180000 40520 6 dmem_dina[24]
port 82 nsew signal output
rlabel metal3 s 179200 41896 180000 42016 6 dmem_dina[25]
port 83 nsew signal output
rlabel metal3 s 179200 43392 180000 43512 6 dmem_dina[26]
port 84 nsew signal output
rlabel metal3 s 179200 44888 180000 45008 6 dmem_dina[27]
port 85 nsew signal output
rlabel metal3 s 179200 46384 180000 46504 6 dmem_dina[28]
port 86 nsew signal output
rlabel metal3 s 179200 47880 180000 48000 6 dmem_dina[29]
port 87 nsew signal output
rlabel metal3 s 179200 7488 180000 7608 6 dmem_dina[2]
port 88 nsew signal output
rlabel metal3 s 179200 49376 180000 49496 6 dmem_dina[30]
port 89 nsew signal output
rlabel metal3 s 179200 50872 180000 50992 6 dmem_dina[31]
port 90 nsew signal output
rlabel metal3 s 179200 8984 180000 9104 6 dmem_dina[3]
port 91 nsew signal output
rlabel metal3 s 179200 10480 180000 10600 6 dmem_dina[4]
port 92 nsew signal output
rlabel metal3 s 179200 11976 180000 12096 6 dmem_dina[5]
port 93 nsew signal output
rlabel metal3 s 179200 13472 180000 13592 6 dmem_dina[6]
port 94 nsew signal output
rlabel metal3 s 179200 14968 180000 15088 6 dmem_dina[7]
port 95 nsew signal output
rlabel metal3 s 179200 16464 180000 16584 6 dmem_dina[8]
port 96 nsew signal output
rlabel metal3 s 179200 17960 180000 18080 6 dmem_dina[9]
port 97 nsew signal output
rlabel metal3 s 179200 52368 180000 52488 6 dmem_dinb[0]
port 98 nsew signal output
rlabel metal3 s 179200 67328 180000 67448 6 dmem_dinb[10]
port 99 nsew signal output
rlabel metal3 s 179200 68824 180000 68944 6 dmem_dinb[11]
port 100 nsew signal output
rlabel metal3 s 179200 70320 180000 70440 6 dmem_dinb[12]
port 101 nsew signal output
rlabel metal3 s 179200 71816 180000 71936 6 dmem_dinb[13]
port 102 nsew signal output
rlabel metal3 s 179200 73312 180000 73432 6 dmem_dinb[14]
port 103 nsew signal output
rlabel metal3 s 179200 74808 180000 74928 6 dmem_dinb[15]
port 104 nsew signal output
rlabel metal3 s 179200 76304 180000 76424 6 dmem_dinb[16]
port 105 nsew signal output
rlabel metal3 s 179200 77800 180000 77920 6 dmem_dinb[17]
port 106 nsew signal output
rlabel metal3 s 179200 79296 180000 79416 6 dmem_dinb[18]
port 107 nsew signal output
rlabel metal3 s 179200 80792 180000 80912 6 dmem_dinb[19]
port 108 nsew signal output
rlabel metal3 s 179200 53864 180000 53984 6 dmem_dinb[1]
port 109 nsew signal output
rlabel metal3 s 179200 82288 180000 82408 6 dmem_dinb[20]
port 110 nsew signal output
rlabel metal3 s 179200 83784 180000 83904 6 dmem_dinb[21]
port 111 nsew signal output
rlabel metal3 s 179200 85280 180000 85400 6 dmem_dinb[22]
port 112 nsew signal output
rlabel metal3 s 179200 86776 180000 86896 6 dmem_dinb[23]
port 113 nsew signal output
rlabel metal3 s 179200 88272 180000 88392 6 dmem_dinb[24]
port 114 nsew signal output
rlabel metal3 s 179200 89768 180000 89888 6 dmem_dinb[25]
port 115 nsew signal output
rlabel metal3 s 179200 91264 180000 91384 6 dmem_dinb[26]
port 116 nsew signal output
rlabel metal3 s 179200 92760 180000 92880 6 dmem_dinb[27]
port 117 nsew signal output
rlabel metal3 s 179200 94256 180000 94376 6 dmem_dinb[28]
port 118 nsew signal output
rlabel metal3 s 179200 95752 180000 95872 6 dmem_dinb[29]
port 119 nsew signal output
rlabel metal3 s 179200 55360 180000 55480 6 dmem_dinb[2]
port 120 nsew signal output
rlabel metal3 s 179200 97248 180000 97368 6 dmem_dinb[30]
port 121 nsew signal output
rlabel metal3 s 179200 98744 180000 98864 6 dmem_dinb[31]
port 122 nsew signal output
rlabel metal3 s 179200 56856 180000 56976 6 dmem_dinb[3]
port 123 nsew signal output
rlabel metal3 s 179200 58352 180000 58472 6 dmem_dinb[4]
port 124 nsew signal output
rlabel metal3 s 179200 59848 180000 59968 6 dmem_dinb[5]
port 125 nsew signal output
rlabel metal3 s 179200 61344 180000 61464 6 dmem_dinb[6]
port 126 nsew signal output
rlabel metal3 s 179200 62840 180000 62960 6 dmem_dinb[7]
port 127 nsew signal output
rlabel metal3 s 179200 64336 180000 64456 6 dmem_dinb[8]
port 128 nsew signal output
rlabel metal3 s 179200 65832 180000 65952 6 dmem_dinb[9]
port 129 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 dmem_doutb[0]
port 130 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 dmem_doutb[10]
port 131 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 dmem_doutb[11]
port 132 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 dmem_doutb[12]
port 133 nsew signal input
rlabel metal3 s 0 54816 800 54936 6 dmem_doutb[13]
port 134 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 dmem_doutb[14]
port 135 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 dmem_doutb[15]
port 136 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 dmem_doutb[16]
port 137 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 dmem_doutb[17]
port 138 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 dmem_doutb[18]
port 139 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 dmem_doutb[19]
port 140 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 dmem_doutb[1]
port 141 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 dmem_doutb[20]
port 142 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 dmem_doutb[21]
port 143 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 dmem_doutb[22]
port 144 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 dmem_doutb[23]
port 145 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 dmem_doutb[24]
port 146 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 dmem_doutb[25]
port 147 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 dmem_doutb[26]
port 148 nsew signal input
rlabel metal3 s 0 102416 800 102536 6 dmem_doutb[27]
port 149 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 dmem_doutb[28]
port 150 nsew signal input
rlabel metal3 s 0 109216 800 109336 6 dmem_doutb[29]
port 151 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 dmem_doutb[2]
port 152 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 dmem_doutb[30]
port 153 nsew signal input
rlabel metal3 s 0 116016 800 116136 6 dmem_doutb[31]
port 154 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 dmem_doutb[3]
port 155 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 dmem_doutb[4]
port 156 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 dmem_doutb[5]
port 157 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 dmem_doutb[6]
port 158 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 dmem_doutb[7]
port 159 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 dmem_doutb[8]
port 160 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 dmem_doutb[9]
port 161 nsew signal input
rlabel metal3 s 179200 113704 180000 113824 6 dmem_ena
port 162 nsew signal output
rlabel metal3 s 179200 115200 180000 115320 6 dmem_enb
port 163 nsew signal output
rlabel metal3 s 179200 100240 180000 100360 6 dmem_wea0
port 164 nsew signal output
rlabel metal3 s 179200 101736 180000 101856 6 dmem_wea[0]
port 165 nsew signal output
rlabel metal3 s 179200 104728 180000 104848 6 dmem_wea[1]
port 166 nsew signal output
rlabel metal3 s 179200 107720 180000 107840 6 dmem_wea[2]
port 167 nsew signal output
rlabel metal3 s 179200 110712 180000 110832 6 dmem_wea[3]
port 168 nsew signal output
rlabel metal3 s 179200 103232 180000 103352 6 dmem_web[0]
port 169 nsew signal output
rlabel metal3 s 179200 106224 180000 106344 6 dmem_web[1]
port 170 nsew signal output
rlabel metal3 s 179200 109216 180000 109336 6 dmem_web[2]
port 171 nsew signal output
rlabel metal3 s 179200 112208 180000 112328 6 dmem_web[3]
port 172 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 imem_addr[0]
port 173 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 imem_addr[10]
port 174 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 imem_addr[11]
port 175 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 imem_addr[12]
port 176 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 imem_addr[13]
port 177 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 imem_addr[14]
port 178 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 imem_addr[15]
port 179 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 imem_addr[16]
port 180 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 imem_addr[17]
port 181 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 imem_addr[18]
port 182 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 imem_addr[19]
port 183 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 imem_addr[1]
port 184 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 imem_addr[20]
port 185 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 imem_addr[21]
port 186 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 imem_addr[22]
port 187 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 imem_addr[23]
port 188 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 imem_addr[24]
port 189 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 imem_addr[25]
port 190 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 imem_addr[26]
port 191 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 imem_addr[27]
port 192 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 imem_addr[28]
port 193 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 imem_addr[29]
port 194 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 imem_addr[2]
port 195 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 imem_addr[30]
port 196 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 imem_addr[31]
port 197 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 imem_addr[3]
port 198 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 imem_addr[4]
port 199 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 imem_addr[5]
port 200 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 imem_addr[6]
port 201 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 imem_addr[7]
port 202 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 imem_addr[8]
port 203 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 imem_addr[9]
port 204 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 imem_data[0]
port 205 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 imem_data[10]
port 206 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 imem_data[11]
port 207 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 imem_data[12]
port 208 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 imem_data[13]
port 209 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 imem_data[14]
port 210 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 imem_data[15]
port 211 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 imem_data[16]
port 212 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 imem_data[17]
port 213 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 imem_data[18]
port 214 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 imem_data[19]
port 215 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 imem_data[1]
port 216 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 imem_data[20]
port 217 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 imem_data[21]
port 218 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 imem_data[22]
port 219 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 imem_data[23]
port 220 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 imem_data[24]
port 221 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 imem_data[25]
port 222 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 imem_data[26]
port 223 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 imem_data[27]
port 224 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 imem_data[28]
port 225 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 imem_data[29]
port 226 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 imem_data[2]
port 227 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 imem_data[30]
port 228 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 imem_data[31]
port 229 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 imem_data[3]
port 230 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 imem_data[4]
port 231 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 imem_data[5]
port 232 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 imem_data[6]
port 233 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 imem_data[7]
port 234 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 imem_data[8]
port 235 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 imem_data[9]
port 236 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 reset
port 237 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 238 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 238 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 238 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 238 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 238 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 238 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 239 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 239 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 239 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 239 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 239 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 239 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 48766322
string GDS_FILE /home/ali11-2000/efabless/mpw-waprv/openlane/warpv_core/runs/22_09_11_16_35/results/signoff/warpv_core.magic.gds
string GDS_START 1305772
<< end >>

