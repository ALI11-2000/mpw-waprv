VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_interface
  CLASS BLOCK ;
  FOREIGN wb_interface ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 397.160 500.000 397.760 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 406.680 500.000 407.280 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 416.200 500.000 416.800 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 425.720 500.000 426.320 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 435.240 500.000 435.840 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 444.760 500.000 445.360 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 454.280 500.000 454.880 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 463.800 500.000 464.400 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 473.320 500.000 473.920 ;
    END
  END addr0[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 25.880 500.000 26.480 ;
    END
  END clk0
  PIN csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 35.400 500.000 36.000 ;
    END
  END csb0
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 92.520 500.000 93.120 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.720 500.000 188.320 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 197.240 500.000 197.840 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 206.760 500.000 207.360 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 216.280 500.000 216.880 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 225.800 500.000 226.400 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 235.320 500.000 235.920 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 244.840 500.000 245.440 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 254.360 500.000 254.960 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 263.880 500.000 264.480 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 273.400 500.000 274.000 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.040 500.000 102.640 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 282.920 500.000 283.520 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 292.440 500.000 293.040 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 301.960 500.000 302.560 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 311.480 500.000 312.080 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 321.000 500.000 321.600 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 330.520 500.000 331.120 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 349.560 500.000 350.160 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 359.080 500.000 359.680 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 368.600 500.000 369.200 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 111.560 500.000 112.160 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 378.120 500.000 378.720 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 387.640 500.000 388.240 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 121.080 500.000 121.680 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 130.600 500.000 131.200 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 140.120 500.000 140.720 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 149.640 500.000 150.240 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 159.160 500.000 159.760 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 168.680 500.000 169.280 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 178.200 500.000 178.800 ;
    END
  END din0[9]
  PIN dmem_addrb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 496.000 17.390 500.000 ;
    END
  END dmem_addrb[0]
  PIN dmem_addrb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 496.000 47.750 500.000 ;
    END
  END dmem_addrb[1]
  PIN dmem_addrb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 496.000 78.110 500.000 ;
    END
  END dmem_addrb[2]
  PIN dmem_addrb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 496.000 108.470 500.000 ;
    END
  END dmem_addrb[3]
  PIN dmem_addrb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 496.000 138.830 500.000 ;
    END
  END dmem_addrb[4]
  PIN dmem_addrb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 496.000 169.190 500.000 ;
    END
  END dmem_addrb[5]
  PIN dmem_addrb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 496.000 199.550 500.000 ;
    END
  END dmem_addrb[6]
  PIN dmem_addrb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 496.000 229.910 500.000 ;
    END
  END dmem_addrb[7]
  PIN dmem_addrb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 496.000 27.510 500.000 ;
    END
  END dmem_addrb_o[0]
  PIN dmem_addrb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 496.000 57.870 500.000 ;
    END
  END dmem_addrb_o[1]
  PIN dmem_addrb_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 496.000 88.230 500.000 ;
    END
  END dmem_addrb_o[2]
  PIN dmem_addrb_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 496.000 118.590 500.000 ;
    END
  END dmem_addrb_o[3]
  PIN dmem_addrb_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 496.000 148.950 500.000 ;
    END
  END dmem_addrb_o[4]
  PIN dmem_addrb_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 496.000 179.310 500.000 ;
    END
  END dmem_addrb_o[5]
  PIN dmem_addrb_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 496.000 209.670 500.000 ;
    END
  END dmem_addrb_o[6]
  PIN dmem_addrb_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 496.000 240.030 500.000 ;
    END
  END dmem_addrb_o[7]
  PIN dmem_doutb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 496.000 37.630 500.000 ;
    END
  END dmem_doutb[0]
  PIN dmem_doutb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 496.000 280.510 500.000 ;
    END
  END dmem_doutb[10]
  PIN dmem_doutb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 496.000 290.630 500.000 ;
    END
  END dmem_doutb[11]
  PIN dmem_doutb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 496.000 300.750 500.000 ;
    END
  END dmem_doutb[12]
  PIN dmem_doutb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 496.000 310.870 500.000 ;
    END
  END dmem_doutb[13]
  PIN dmem_doutb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 496.000 320.990 500.000 ;
    END
  END dmem_doutb[14]
  PIN dmem_doutb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 496.000 331.110 500.000 ;
    END
  END dmem_doutb[15]
  PIN dmem_doutb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 496.000 341.230 500.000 ;
    END
  END dmem_doutb[16]
  PIN dmem_doutb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 496.000 351.350 500.000 ;
    END
  END dmem_doutb[17]
  PIN dmem_doutb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 496.000 361.470 500.000 ;
    END
  END dmem_doutb[18]
  PIN dmem_doutb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 496.000 371.590 500.000 ;
    END
  END dmem_doutb[19]
  PIN dmem_doutb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 496.000 67.990 500.000 ;
    END
  END dmem_doutb[1]
  PIN dmem_doutb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 496.000 381.710 500.000 ;
    END
  END dmem_doutb[20]
  PIN dmem_doutb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 496.000 391.830 500.000 ;
    END
  END dmem_doutb[21]
  PIN dmem_doutb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 496.000 401.950 500.000 ;
    END
  END dmem_doutb[22]
  PIN dmem_doutb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 496.000 412.070 500.000 ;
    END
  END dmem_doutb[23]
  PIN dmem_doutb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 496.000 422.190 500.000 ;
    END
  END dmem_doutb[24]
  PIN dmem_doutb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 496.000 432.310 500.000 ;
    END
  END dmem_doutb[25]
  PIN dmem_doutb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 496.000 442.430 500.000 ;
    END
  END dmem_doutb[26]
  PIN dmem_doutb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 496.000 452.550 500.000 ;
    END
  END dmem_doutb[27]
  PIN dmem_doutb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 496.000 462.670 500.000 ;
    END
  END dmem_doutb[28]
  PIN dmem_doutb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 496.000 472.790 500.000 ;
    END
  END dmem_doutb[29]
  PIN dmem_doutb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 496.000 98.350 500.000 ;
    END
  END dmem_doutb[2]
  PIN dmem_doutb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 496.000 482.910 500.000 ;
    END
  END dmem_doutb[30]
  PIN dmem_doutb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 496.000 493.030 500.000 ;
    END
  END dmem_doutb[31]
  PIN dmem_doutb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 496.000 128.710 500.000 ;
    END
  END dmem_doutb[3]
  PIN dmem_doutb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 496.000 159.070 500.000 ;
    END
  END dmem_doutb[4]
  PIN dmem_doutb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 496.000 189.430 500.000 ;
    END
  END dmem_doutb[5]
  PIN dmem_doutb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 496.000 219.790 500.000 ;
    END
  END dmem_doutb[6]
  PIN dmem_doutb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 496.000 250.150 500.000 ;
    END
  END dmem_doutb[7]
  PIN dmem_doutb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 496.000 260.270 500.000 ;
    END
  END dmem_doutb[8]
  PIN dmem_doutb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 496.000 270.390 500.000 ;
    END
  END dmem_doutb[9]
  PIN dmem_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 496.000 7.270 500.000 ;
    END
  END dmem_enb
  PIN imem_rd_cs1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 16.360 500.000 16.960 ;
    END
  END imem_rd_cs1
  PIN processor_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 482.840 500.000 483.440 ;
    END
  END processor_reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END wbs_we_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.920 500.000 45.520 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 54.440 500.000 55.040 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 63.960 500.000 64.560 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 73.480 500.000 74.080 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 83.000 500.000 83.600 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 7.550 495.720 16.830 496.810 ;
        RECT 17.670 495.720 26.950 496.810 ;
        RECT 27.790 495.720 37.070 496.810 ;
        RECT 37.910 495.720 47.190 496.810 ;
        RECT 48.030 495.720 57.310 496.810 ;
        RECT 58.150 495.720 67.430 496.810 ;
        RECT 68.270 495.720 77.550 496.810 ;
        RECT 78.390 495.720 87.670 496.810 ;
        RECT 88.510 495.720 97.790 496.810 ;
        RECT 98.630 495.720 107.910 496.810 ;
        RECT 108.750 495.720 118.030 496.810 ;
        RECT 118.870 495.720 128.150 496.810 ;
        RECT 128.990 495.720 138.270 496.810 ;
        RECT 139.110 495.720 148.390 496.810 ;
        RECT 149.230 495.720 158.510 496.810 ;
        RECT 159.350 495.720 168.630 496.810 ;
        RECT 169.470 495.720 178.750 496.810 ;
        RECT 179.590 495.720 188.870 496.810 ;
        RECT 189.710 495.720 198.990 496.810 ;
        RECT 199.830 495.720 209.110 496.810 ;
        RECT 209.950 495.720 219.230 496.810 ;
        RECT 220.070 495.720 229.350 496.810 ;
        RECT 230.190 495.720 239.470 496.810 ;
        RECT 240.310 495.720 249.590 496.810 ;
        RECT 250.430 495.720 259.710 496.810 ;
        RECT 260.550 495.720 269.830 496.810 ;
        RECT 270.670 495.720 279.950 496.810 ;
        RECT 280.790 495.720 290.070 496.810 ;
        RECT 290.910 495.720 300.190 496.810 ;
        RECT 301.030 495.720 310.310 496.810 ;
        RECT 311.150 495.720 320.430 496.810 ;
        RECT 321.270 495.720 330.550 496.810 ;
        RECT 331.390 495.720 340.670 496.810 ;
        RECT 341.510 495.720 350.790 496.810 ;
        RECT 351.630 495.720 360.910 496.810 ;
        RECT 361.750 495.720 371.030 496.810 ;
        RECT 371.870 495.720 381.150 496.810 ;
        RECT 381.990 495.720 391.270 496.810 ;
        RECT 392.110 495.720 401.390 496.810 ;
        RECT 402.230 495.720 411.510 496.810 ;
        RECT 412.350 495.720 421.630 496.810 ;
        RECT 422.470 495.720 431.750 496.810 ;
        RECT 432.590 495.720 441.870 496.810 ;
        RECT 442.710 495.720 451.990 496.810 ;
        RECT 452.830 495.720 462.110 496.810 ;
        RECT 462.950 495.720 472.230 496.810 ;
        RECT 473.070 495.720 482.350 496.810 ;
        RECT 483.190 495.720 492.470 496.810 ;
        RECT 6.990 10.695 493.020 495.720 ;
      LAYER met3 ;
        RECT 4.000 483.840 496.000 487.045 ;
        RECT 4.000 482.440 495.600 483.840 ;
        RECT 4.000 474.320 496.000 482.440 ;
        RECT 4.000 472.920 495.600 474.320 ;
        RECT 4.000 464.800 496.000 472.920 ;
        RECT 4.400 463.400 495.600 464.800 ;
        RECT 4.000 460.720 496.000 463.400 ;
        RECT 4.400 459.320 496.000 460.720 ;
        RECT 4.000 456.640 496.000 459.320 ;
        RECT 4.400 455.280 496.000 456.640 ;
        RECT 4.400 455.240 495.600 455.280 ;
        RECT 4.000 453.880 495.600 455.240 ;
        RECT 4.000 452.560 496.000 453.880 ;
        RECT 4.400 451.160 496.000 452.560 ;
        RECT 4.000 448.480 496.000 451.160 ;
        RECT 4.400 447.080 496.000 448.480 ;
        RECT 4.000 445.760 496.000 447.080 ;
        RECT 4.000 444.400 495.600 445.760 ;
        RECT 4.400 444.360 495.600 444.400 ;
        RECT 4.400 443.000 496.000 444.360 ;
        RECT 4.000 440.320 496.000 443.000 ;
        RECT 4.400 438.920 496.000 440.320 ;
        RECT 4.000 436.240 496.000 438.920 ;
        RECT 4.400 434.840 495.600 436.240 ;
        RECT 4.000 432.160 496.000 434.840 ;
        RECT 4.400 430.760 496.000 432.160 ;
        RECT 4.000 428.080 496.000 430.760 ;
        RECT 4.400 426.720 496.000 428.080 ;
        RECT 4.400 426.680 495.600 426.720 ;
        RECT 4.000 425.320 495.600 426.680 ;
        RECT 4.000 424.000 496.000 425.320 ;
        RECT 4.400 422.600 496.000 424.000 ;
        RECT 4.000 419.920 496.000 422.600 ;
        RECT 4.400 418.520 496.000 419.920 ;
        RECT 4.000 417.200 496.000 418.520 ;
        RECT 4.000 415.840 495.600 417.200 ;
        RECT 4.400 415.800 495.600 415.840 ;
        RECT 4.400 414.440 496.000 415.800 ;
        RECT 4.000 411.760 496.000 414.440 ;
        RECT 4.400 410.360 496.000 411.760 ;
        RECT 4.000 407.680 496.000 410.360 ;
        RECT 4.400 406.280 495.600 407.680 ;
        RECT 4.000 403.600 496.000 406.280 ;
        RECT 4.400 402.200 496.000 403.600 ;
        RECT 4.000 399.520 496.000 402.200 ;
        RECT 4.400 398.160 496.000 399.520 ;
        RECT 4.400 398.120 495.600 398.160 ;
        RECT 4.000 396.760 495.600 398.120 ;
        RECT 4.000 395.440 496.000 396.760 ;
        RECT 4.400 394.040 496.000 395.440 ;
        RECT 4.000 391.360 496.000 394.040 ;
        RECT 4.400 389.960 496.000 391.360 ;
        RECT 4.000 388.640 496.000 389.960 ;
        RECT 4.000 387.280 495.600 388.640 ;
        RECT 4.400 387.240 495.600 387.280 ;
        RECT 4.400 385.880 496.000 387.240 ;
        RECT 4.000 383.200 496.000 385.880 ;
        RECT 4.400 381.800 496.000 383.200 ;
        RECT 4.000 379.120 496.000 381.800 ;
        RECT 4.400 377.720 495.600 379.120 ;
        RECT 4.000 375.040 496.000 377.720 ;
        RECT 4.400 373.640 496.000 375.040 ;
        RECT 4.000 370.960 496.000 373.640 ;
        RECT 4.400 369.600 496.000 370.960 ;
        RECT 4.400 369.560 495.600 369.600 ;
        RECT 4.000 368.200 495.600 369.560 ;
        RECT 4.000 366.880 496.000 368.200 ;
        RECT 4.400 365.480 496.000 366.880 ;
        RECT 4.000 362.800 496.000 365.480 ;
        RECT 4.400 361.400 496.000 362.800 ;
        RECT 4.000 360.080 496.000 361.400 ;
        RECT 4.000 358.720 495.600 360.080 ;
        RECT 4.400 358.680 495.600 358.720 ;
        RECT 4.400 357.320 496.000 358.680 ;
        RECT 4.000 354.640 496.000 357.320 ;
        RECT 4.400 353.240 496.000 354.640 ;
        RECT 4.000 350.560 496.000 353.240 ;
        RECT 4.400 349.160 495.600 350.560 ;
        RECT 4.000 346.480 496.000 349.160 ;
        RECT 4.400 345.080 496.000 346.480 ;
        RECT 4.000 342.400 496.000 345.080 ;
        RECT 4.400 341.040 496.000 342.400 ;
        RECT 4.400 341.000 495.600 341.040 ;
        RECT 4.000 339.640 495.600 341.000 ;
        RECT 4.000 338.320 496.000 339.640 ;
        RECT 4.400 336.920 496.000 338.320 ;
        RECT 4.000 334.240 496.000 336.920 ;
        RECT 4.400 332.840 496.000 334.240 ;
        RECT 4.000 331.520 496.000 332.840 ;
        RECT 4.000 330.160 495.600 331.520 ;
        RECT 4.400 330.120 495.600 330.160 ;
        RECT 4.400 328.760 496.000 330.120 ;
        RECT 4.000 326.080 496.000 328.760 ;
        RECT 4.400 324.680 496.000 326.080 ;
        RECT 4.000 322.000 496.000 324.680 ;
        RECT 4.400 320.600 495.600 322.000 ;
        RECT 4.000 317.920 496.000 320.600 ;
        RECT 4.400 316.520 496.000 317.920 ;
        RECT 4.000 313.840 496.000 316.520 ;
        RECT 4.400 312.480 496.000 313.840 ;
        RECT 4.400 312.440 495.600 312.480 ;
        RECT 4.000 311.080 495.600 312.440 ;
        RECT 4.000 309.760 496.000 311.080 ;
        RECT 4.400 308.360 496.000 309.760 ;
        RECT 4.000 305.680 496.000 308.360 ;
        RECT 4.400 304.280 496.000 305.680 ;
        RECT 4.000 302.960 496.000 304.280 ;
        RECT 4.000 301.600 495.600 302.960 ;
        RECT 4.400 301.560 495.600 301.600 ;
        RECT 4.400 300.200 496.000 301.560 ;
        RECT 4.000 297.520 496.000 300.200 ;
        RECT 4.400 296.120 496.000 297.520 ;
        RECT 4.000 293.440 496.000 296.120 ;
        RECT 4.400 292.040 495.600 293.440 ;
        RECT 4.000 289.360 496.000 292.040 ;
        RECT 4.400 287.960 496.000 289.360 ;
        RECT 4.000 285.280 496.000 287.960 ;
        RECT 4.400 283.920 496.000 285.280 ;
        RECT 4.400 283.880 495.600 283.920 ;
        RECT 4.000 282.520 495.600 283.880 ;
        RECT 4.000 281.200 496.000 282.520 ;
        RECT 4.400 279.800 496.000 281.200 ;
        RECT 4.000 277.120 496.000 279.800 ;
        RECT 4.400 275.720 496.000 277.120 ;
        RECT 4.000 274.400 496.000 275.720 ;
        RECT 4.000 273.040 495.600 274.400 ;
        RECT 4.400 273.000 495.600 273.040 ;
        RECT 4.400 271.640 496.000 273.000 ;
        RECT 4.000 268.960 496.000 271.640 ;
        RECT 4.400 267.560 496.000 268.960 ;
        RECT 4.000 264.880 496.000 267.560 ;
        RECT 4.400 263.480 495.600 264.880 ;
        RECT 4.000 260.800 496.000 263.480 ;
        RECT 4.400 259.400 496.000 260.800 ;
        RECT 4.000 256.720 496.000 259.400 ;
        RECT 4.400 255.360 496.000 256.720 ;
        RECT 4.400 255.320 495.600 255.360 ;
        RECT 4.000 253.960 495.600 255.320 ;
        RECT 4.000 252.640 496.000 253.960 ;
        RECT 4.400 251.240 496.000 252.640 ;
        RECT 4.000 248.560 496.000 251.240 ;
        RECT 4.400 247.160 496.000 248.560 ;
        RECT 4.000 245.840 496.000 247.160 ;
        RECT 4.000 244.480 495.600 245.840 ;
        RECT 4.400 244.440 495.600 244.480 ;
        RECT 4.400 243.080 496.000 244.440 ;
        RECT 4.000 240.400 496.000 243.080 ;
        RECT 4.400 239.000 496.000 240.400 ;
        RECT 4.000 236.320 496.000 239.000 ;
        RECT 4.400 234.920 495.600 236.320 ;
        RECT 4.000 232.240 496.000 234.920 ;
        RECT 4.400 230.840 496.000 232.240 ;
        RECT 4.000 228.160 496.000 230.840 ;
        RECT 4.400 226.800 496.000 228.160 ;
        RECT 4.400 226.760 495.600 226.800 ;
        RECT 4.000 225.400 495.600 226.760 ;
        RECT 4.000 224.080 496.000 225.400 ;
        RECT 4.400 222.680 496.000 224.080 ;
        RECT 4.000 220.000 496.000 222.680 ;
        RECT 4.400 218.600 496.000 220.000 ;
        RECT 4.000 217.280 496.000 218.600 ;
        RECT 4.000 215.920 495.600 217.280 ;
        RECT 4.400 215.880 495.600 215.920 ;
        RECT 4.400 214.520 496.000 215.880 ;
        RECT 4.000 211.840 496.000 214.520 ;
        RECT 4.400 210.440 496.000 211.840 ;
        RECT 4.000 207.760 496.000 210.440 ;
        RECT 4.400 206.360 495.600 207.760 ;
        RECT 4.000 203.680 496.000 206.360 ;
        RECT 4.400 202.280 496.000 203.680 ;
        RECT 4.000 199.600 496.000 202.280 ;
        RECT 4.400 198.240 496.000 199.600 ;
        RECT 4.400 198.200 495.600 198.240 ;
        RECT 4.000 196.840 495.600 198.200 ;
        RECT 4.000 195.520 496.000 196.840 ;
        RECT 4.400 194.120 496.000 195.520 ;
        RECT 4.000 191.440 496.000 194.120 ;
        RECT 4.400 190.040 496.000 191.440 ;
        RECT 4.000 188.720 496.000 190.040 ;
        RECT 4.000 187.360 495.600 188.720 ;
        RECT 4.400 187.320 495.600 187.360 ;
        RECT 4.400 185.960 496.000 187.320 ;
        RECT 4.000 183.280 496.000 185.960 ;
        RECT 4.400 181.880 496.000 183.280 ;
        RECT 4.000 179.200 496.000 181.880 ;
        RECT 4.400 177.800 495.600 179.200 ;
        RECT 4.000 175.120 496.000 177.800 ;
        RECT 4.400 173.720 496.000 175.120 ;
        RECT 4.000 171.040 496.000 173.720 ;
        RECT 4.400 169.680 496.000 171.040 ;
        RECT 4.400 169.640 495.600 169.680 ;
        RECT 4.000 168.280 495.600 169.640 ;
        RECT 4.000 166.960 496.000 168.280 ;
        RECT 4.400 165.560 496.000 166.960 ;
        RECT 4.000 162.880 496.000 165.560 ;
        RECT 4.400 161.480 496.000 162.880 ;
        RECT 4.000 160.160 496.000 161.480 ;
        RECT 4.000 158.800 495.600 160.160 ;
        RECT 4.400 158.760 495.600 158.800 ;
        RECT 4.400 157.400 496.000 158.760 ;
        RECT 4.000 154.720 496.000 157.400 ;
        RECT 4.400 153.320 496.000 154.720 ;
        RECT 4.000 150.640 496.000 153.320 ;
        RECT 4.400 149.240 495.600 150.640 ;
        RECT 4.000 146.560 496.000 149.240 ;
        RECT 4.400 145.160 496.000 146.560 ;
        RECT 4.000 142.480 496.000 145.160 ;
        RECT 4.400 141.120 496.000 142.480 ;
        RECT 4.400 141.080 495.600 141.120 ;
        RECT 4.000 139.720 495.600 141.080 ;
        RECT 4.000 138.400 496.000 139.720 ;
        RECT 4.400 137.000 496.000 138.400 ;
        RECT 4.000 134.320 496.000 137.000 ;
        RECT 4.400 132.920 496.000 134.320 ;
        RECT 4.000 131.600 496.000 132.920 ;
        RECT 4.000 130.240 495.600 131.600 ;
        RECT 4.400 130.200 495.600 130.240 ;
        RECT 4.400 128.840 496.000 130.200 ;
        RECT 4.000 126.160 496.000 128.840 ;
        RECT 4.400 124.760 496.000 126.160 ;
        RECT 4.000 122.080 496.000 124.760 ;
        RECT 4.400 120.680 495.600 122.080 ;
        RECT 4.000 118.000 496.000 120.680 ;
        RECT 4.400 116.600 496.000 118.000 ;
        RECT 4.000 113.920 496.000 116.600 ;
        RECT 4.400 112.560 496.000 113.920 ;
        RECT 4.400 112.520 495.600 112.560 ;
        RECT 4.000 111.160 495.600 112.520 ;
        RECT 4.000 109.840 496.000 111.160 ;
        RECT 4.400 108.440 496.000 109.840 ;
        RECT 4.000 105.760 496.000 108.440 ;
        RECT 4.400 104.360 496.000 105.760 ;
        RECT 4.000 103.040 496.000 104.360 ;
        RECT 4.000 101.680 495.600 103.040 ;
        RECT 4.400 101.640 495.600 101.680 ;
        RECT 4.400 100.280 496.000 101.640 ;
        RECT 4.000 97.600 496.000 100.280 ;
        RECT 4.400 96.200 496.000 97.600 ;
        RECT 4.000 93.520 496.000 96.200 ;
        RECT 4.400 92.120 495.600 93.520 ;
        RECT 4.000 89.440 496.000 92.120 ;
        RECT 4.400 88.040 496.000 89.440 ;
        RECT 4.000 85.360 496.000 88.040 ;
        RECT 4.400 84.000 496.000 85.360 ;
        RECT 4.400 83.960 495.600 84.000 ;
        RECT 4.000 82.600 495.600 83.960 ;
        RECT 4.000 81.280 496.000 82.600 ;
        RECT 4.400 79.880 496.000 81.280 ;
        RECT 4.000 77.200 496.000 79.880 ;
        RECT 4.400 75.800 496.000 77.200 ;
        RECT 4.000 74.480 496.000 75.800 ;
        RECT 4.000 73.120 495.600 74.480 ;
        RECT 4.400 73.080 495.600 73.120 ;
        RECT 4.400 71.720 496.000 73.080 ;
        RECT 4.000 69.040 496.000 71.720 ;
        RECT 4.400 67.640 496.000 69.040 ;
        RECT 4.000 64.960 496.000 67.640 ;
        RECT 4.400 63.560 495.600 64.960 ;
        RECT 4.000 60.880 496.000 63.560 ;
        RECT 4.400 59.480 496.000 60.880 ;
        RECT 4.000 56.800 496.000 59.480 ;
        RECT 4.400 55.440 496.000 56.800 ;
        RECT 4.400 55.400 495.600 55.440 ;
        RECT 4.000 54.040 495.600 55.400 ;
        RECT 4.000 52.720 496.000 54.040 ;
        RECT 4.400 51.320 496.000 52.720 ;
        RECT 4.000 48.640 496.000 51.320 ;
        RECT 4.400 47.240 496.000 48.640 ;
        RECT 4.000 45.920 496.000 47.240 ;
        RECT 4.000 44.560 495.600 45.920 ;
        RECT 4.400 44.520 495.600 44.560 ;
        RECT 4.400 43.160 496.000 44.520 ;
        RECT 4.000 40.480 496.000 43.160 ;
        RECT 4.400 39.080 496.000 40.480 ;
        RECT 4.000 36.400 496.000 39.080 ;
        RECT 4.400 35.000 495.600 36.400 ;
        RECT 4.000 26.880 496.000 35.000 ;
        RECT 4.000 25.480 495.600 26.880 ;
        RECT 4.000 17.360 496.000 25.480 ;
        RECT 4.000 15.960 495.600 17.360 ;
        RECT 4.000 10.715 496.000 15.960 ;
  END
END wb_interface
END LIBRARY

