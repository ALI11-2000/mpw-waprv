* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for wb_interface abstract view
.subckt wb_interface addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] addr0[8] clk0 csb0 din0[0] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[1] din0[20] din0[21] din0[22]
+ din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[2] din0[30]
+ din0[31] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] imem_rd_cs1 processor_reset
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i web0 wmask0[0]
+ wmask0[1] wmask0[2] wmask0[3]
.ends

* Black-box entry subcircuit for sky130_sram_1kbyte_1rw1r_32x256_8 abstract view
.subckt sky130_sram_1kbyte_1rw1r_32x256_8 din0[0] din0[1] din0[2] din0[3] din0[4]
+ din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr1[0] addr1[1]
+ addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] csb0 csb1 web0 clk0 clk1 wmask0[0]
+ wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5]
+ dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14]
+ dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22]
+ dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30]
+ dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7]
+ dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16]
+ dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24]
+ dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31] vccd1 vssd1
.ends

* Black-box entry subcircuit for warpv_core abstract view
.subckt warpv_core clk dmem_addra[0] dmem_addra[10] dmem_addra[11] dmem_addra[12]
+ dmem_addra[13] dmem_addra[14] dmem_addra[15] dmem_addra[16] dmem_addra[17] dmem_addra[18]
+ dmem_addra[19] dmem_addra[1] dmem_addra[20] dmem_addra[21] dmem_addra[22] dmem_addra[23]
+ dmem_addra[24] dmem_addra[25] dmem_addra[26] dmem_addra[27] dmem_addra[28] dmem_addra[29]
+ dmem_addra[2] dmem_addra[30] dmem_addra[31] dmem_addra[3] dmem_addra[4] dmem_addra[5]
+ dmem_addra[6] dmem_addra[7] dmem_addra[8] dmem_addra[9] dmem_addrb[0] dmem_addrb[10]
+ dmem_addrb[11] dmem_addrb[12] dmem_addrb[13] dmem_addrb[14] dmem_addrb[15] dmem_addrb[16]
+ dmem_addrb[17] dmem_addrb[18] dmem_addrb[19] dmem_addrb[1] dmem_addrb[20] dmem_addrb[21]
+ dmem_addrb[22] dmem_addrb[23] dmem_addrb[24] dmem_addrb[25] dmem_addrb[26] dmem_addrb[27]
+ dmem_addrb[28] dmem_addrb[29] dmem_addrb[2] dmem_addrb[30] dmem_addrb[31] dmem_addrb[3]
+ dmem_addrb[4] dmem_addrb[5] dmem_addrb[6] dmem_addrb[7] dmem_addrb[8] dmem_addrb[9]
+ dmem_dina[0] dmem_dina[10] dmem_dina[11] dmem_dina[12] dmem_dina[13] dmem_dina[14]
+ dmem_dina[15] dmem_dina[16] dmem_dina[17] dmem_dina[18] dmem_dina[19] dmem_dina[1]
+ dmem_dina[20] dmem_dina[21] dmem_dina[22] dmem_dina[23] dmem_dina[24] dmem_dina[25]
+ dmem_dina[26] dmem_dina[27] dmem_dina[28] dmem_dina[29] dmem_dina[2] dmem_dina[30]
+ dmem_dina[31] dmem_dina[3] dmem_dina[4] dmem_dina[5] dmem_dina[6] dmem_dina[7] dmem_dina[8]
+ dmem_dina[9] dmem_dinb[0] dmem_dinb[10] dmem_dinb[11] dmem_dinb[12] dmem_dinb[13]
+ dmem_dinb[14] dmem_dinb[15] dmem_dinb[16] dmem_dinb[17] dmem_dinb[18] dmem_dinb[19]
+ dmem_dinb[1] dmem_dinb[20] dmem_dinb[21] dmem_dinb[22] dmem_dinb[23] dmem_dinb[24]
+ dmem_dinb[25] dmem_dinb[26] dmem_dinb[27] dmem_dinb[28] dmem_dinb[29] dmem_dinb[2]
+ dmem_dinb[30] dmem_dinb[31] dmem_dinb[3] dmem_dinb[4] dmem_dinb[5] dmem_dinb[6]
+ dmem_dinb[7] dmem_dinb[8] dmem_dinb[9] dmem_doutb[0] dmem_doutb[10] dmem_doutb[11]
+ dmem_doutb[12] dmem_doutb[13] dmem_doutb[14] dmem_doutb[15] dmem_doutb[16] dmem_doutb[17]
+ dmem_doutb[18] dmem_doutb[19] dmem_doutb[1] dmem_doutb[20] dmem_doutb[21] dmem_doutb[22]
+ dmem_doutb[23] dmem_doutb[24] dmem_doutb[25] dmem_doutb[26] dmem_doutb[27] dmem_doutb[28]
+ dmem_doutb[29] dmem_doutb[2] dmem_doutb[30] dmem_doutb[31] dmem_doutb[3] dmem_doutb[4]
+ dmem_doutb[5] dmem_doutb[6] dmem_doutb[7] dmem_doutb[8] dmem_doutb[9] dmem_ena dmem_enb
+ dmem_wea0 dmem_wea[0] dmem_wea[1] dmem_wea[2] dmem_wea[3] dmem_web[0] dmem_web[1]
+ dmem_web[2] dmem_web[3] imem_addr[0] imem_addr[10] imem_addr[11] imem_addr[12] imem_addr[13]
+ imem_addr[14] imem_addr[15] imem_addr[16] imem_addr[17] imem_addr[18] imem_addr[19]
+ imem_addr[1] imem_addr[20] imem_addr[21] imem_addr[22] imem_addr[23] imem_addr[24]
+ imem_addr[25] imem_addr[26] imem_addr[27] imem_addr[28] imem_addr[29] imem_addr[2]
+ imem_addr[30] imem_addr[31] imem_addr[3] imem_addr[4] imem_addr[5] imem_addr[6]
+ imem_addr[7] imem_addr[8] imem_addr[9] imem_data[0] imem_data[10] imem_data[11]
+ imem_data[12] imem_data[13] imem_data[14] imem_data[15] imem_data[16] imem_data[17]
+ imem_data[18] imem_data[19] imem_data[1] imem_data[20] imem_data[21] imem_data[22]
+ imem_data[23] imem_data[24] imem_data[25] imem_data[26] imem_data[27] imem_data[28]
+ imem_data[29] imem_data[2] imem_data[30] imem_data[31] imem_data[3] imem_data[4]
+ imem_data[5] imem_data[6] imem_data[7] imem_data[8] imem_data[9] reset vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xwbs_int la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108]
+ la_data_out[109] la_data_out[110] la_data_out[111] wbs_int/addr0[8] wbs_int/clk0
+ imem/csb0 la_data_out[72] la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85]
+ la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[90]
+ la_data_out[91] la_data_out[73] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[100] la_data_out[101] la_data_out[74] la_data_out[102] la_data_out[103]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[80] la_data_out[81] imem/csb1 core/reset vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i imem/web0 imem/wmask0[0] imem/wmask0[1] imem/wmask0[2] imem/wmask0[3]
+ wb_interface
Ximem la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[110] la_data_out[111]
+ imem/addr1[0] imem/addr1[1] imem/addr1[2] imem/addr1[3] imem/addr1[4] imem/addr1[5]
+ imem/addr1[6] imem/addr1[7] imem/csb0 imem/csb1 imem/web0 wb_clk_i wb_clk_i imem/wmask0[0]
+ imem/wmask0[1] imem/wmask0[2] imem/wmask0[3] imem/dout0[0] imem/dout0[1] imem/dout0[2]
+ imem/dout0[3] imem/dout0[4] imem/dout0[5] imem/dout0[6] imem/dout0[7] imem/dout0[8]
+ imem/dout0[9] imem/dout0[10] imem/dout0[11] imem/dout0[12] imem/dout0[13] imem/dout0[14]
+ imem/dout0[15] imem/dout0[16] imem/dout0[17] imem/dout0[18] imem/dout0[19] imem/dout0[20]
+ imem/dout0[21] imem/dout0[22] imem/dout0[23] imem/dout0[24] imem/dout0[25] imem/dout0[26]
+ imem/dout0[27] imem/dout0[28] imem/dout0[29] imem/dout0[30] imem/dout0[31] imem/dout1[0]
+ imem/dout1[1] imem/dout1[2] imem/dout1[3] imem/dout1[4] imem/dout1[5] imem/dout1[6]
+ imem/dout1[7] imem/dout1[8] imem/dout1[9] imem/dout1[10] imem/dout1[11] imem/dout1[12]
+ imem/dout1[13] imem/dout1[14] imem/dout1[15] imem/dout1[16] imem/dout1[17] imem/dout1[18]
+ imem/dout1[19] imem/dout1[20] imem/dout1[21] imem/dout1[22] imem/dout1[23] imem/dout1[24]
+ imem/dout1[25] imem/dout1[26] imem/dout1[27] imem/dout1[28] imem/dout1[29] imem/dout1[30]
+ imem/dout1[31] vccd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xcore wb_clk_i la_data_out[64] core/dmem_addra[10] core/dmem_addra[11] core/dmem_addra[12]
+ core/dmem_addra[13] core/dmem_addra[14] core/dmem_addra[15] core/dmem_addra[16]
+ core/dmem_addra[17] core/dmem_addra[18] core/dmem_addra[19] la_data_out[65] core/dmem_addra[20]
+ core/dmem_addra[21] core/dmem_addra[22] core/dmem_addra[23] core/dmem_addra[24]
+ core/dmem_addra[25] core/dmem_addra[26] core/dmem_addra[27] core/dmem_addra[28]
+ core/dmem_addra[29] la_data_out[66] core/dmem_addra[30] core/dmem_addra[31] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[70] la_data_out[71] core/dmem_addra[8]
+ core/dmem_addra[9] dmem/addr1[0] core/dmem_addrb[10] core/dmem_addrb[11] core/dmem_addrb[12]
+ core/dmem_addrb[13] core/dmem_addrb[14] core/dmem_addrb[15] core/dmem_addrb[16]
+ core/dmem_addrb[17] core/dmem_addrb[18] core/dmem_addrb[19] dmem/addr1[1] core/dmem_addrb[20]
+ core/dmem_addrb[21] core/dmem_addrb[22] core/dmem_addrb[23] core/dmem_addrb[24]
+ core/dmem_addrb[25] core/dmem_addrb[26] core/dmem_addrb[27] core/dmem_addrb[28]
+ core/dmem_addrb[29] dmem/addr1[2] core/dmem_addrb[30] core/dmem_addrb[31] dmem/addr1[3]
+ dmem/addr1[4] dmem/addr1[5] dmem/addr1[6] dmem/addr1[7] core/dmem_addrb[8] core/dmem_addrb[9]
+ la_data_out[32] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[50]
+ la_data_out[51] la_data_out[33] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[60] la_data_out[61] la_data_out[34] la_data_out[62] la_data_out[63]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[40] la_data_out[41] core/dmem_dinb[0] core/dmem_dinb[10] core/dmem_dinb[11]
+ core/dmem_dinb[12] core/dmem_dinb[13] core/dmem_dinb[14] core/dmem_dinb[15] core/dmem_dinb[16]
+ core/dmem_dinb[17] core/dmem_dinb[18] core/dmem_dinb[19] core/dmem_dinb[1] core/dmem_dinb[20]
+ core/dmem_dinb[21] core/dmem_dinb[22] core/dmem_dinb[23] core/dmem_dinb[24] core/dmem_dinb[25]
+ core/dmem_dinb[26] core/dmem_dinb[27] core/dmem_dinb[28] core/dmem_dinb[29] core/dmem_dinb[2]
+ core/dmem_dinb[30] core/dmem_dinb[31] core/dmem_dinb[3] core/dmem_dinb[4] core/dmem_dinb[5]
+ core/dmem_dinb[6] core/dmem_dinb[7] core/dmem_dinb[8] core/dmem_dinb[9] la_data_out[0]
+ la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3] la_data_out[4] la_data_out[5]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] dmem/csb0 dmem/csb1
+ dmem/web0 dmem/wmask0[0] dmem/wmask0[1] dmem/wmask0[2] dmem/wmask0[3] core/dmem_web[0]
+ core/dmem_web[1] core/dmem_web[2] core/dmem_web[3] imem/addr1[0] core/imem_addr[10]
+ core/imem_addr[11] core/imem_addr[12] core/imem_addr[13] core/imem_addr[14] core/imem_addr[15]
+ core/imem_addr[16] core/imem_addr[17] core/imem_addr[18] core/imem_addr[19] imem/addr1[1]
+ core/imem_addr[20] core/imem_addr[21] core/imem_addr[22] core/imem_addr[23] core/imem_addr[24]
+ core/imem_addr[25] core/imem_addr[26] core/imem_addr[27] core/imem_addr[28] core/imem_addr[29]
+ imem/addr1[2] core/imem_addr[30] core/imem_addr[31] imem/addr1[3] imem/addr1[4]
+ imem/addr1[5] imem/addr1[6] imem/addr1[7] core/imem_addr[8] core/imem_addr[9] imem/dout1[0]
+ imem/dout1[10] imem/dout1[11] imem/dout1[12] imem/dout1[13] imem/dout1[14] imem/dout1[15]
+ imem/dout1[16] imem/dout1[17] imem/dout1[18] imem/dout1[19] imem/dout1[1] imem/dout1[20]
+ imem/dout1[21] imem/dout1[22] imem/dout1[23] imem/dout1[24] imem/dout1[25] imem/dout1[26]
+ imem/dout1[27] imem/dout1[28] imem/dout1[29] imem/dout1[2] imem/dout1[30] imem/dout1[31]
+ imem/dout1[3] imem/dout1[4] imem/dout1[5] imem/dout1[6] imem/dout1[7] imem/dout1[8]
+ imem/dout1[9] core/reset vccd1 vssd1 warpv_core
Xdmem la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[70] la_data_out[71]
+ dmem/addr1[0] dmem/addr1[1] dmem/addr1[2] dmem/addr1[3] dmem/addr1[4] dmem/addr1[5]
+ dmem/addr1[6] dmem/addr1[7] dmem/csb0 dmem/csb1 dmem/web0 wb_clk_i wb_clk_i dmem/wmask0[0]
+ dmem/wmask0[1] dmem/wmask0[2] dmem/wmask0[3] dmem/dout0[0] dmem/dout0[1] dmem/dout0[2]
+ dmem/dout0[3] dmem/dout0[4] dmem/dout0[5] dmem/dout0[6] dmem/dout0[7] dmem/dout0[8]
+ dmem/dout0[9] dmem/dout0[10] dmem/dout0[11] dmem/dout0[12] dmem/dout0[13] dmem/dout0[14]
+ dmem/dout0[15] dmem/dout0[16] dmem/dout0[17] dmem/dout0[18] dmem/dout0[19] dmem/dout0[20]
+ dmem/dout0[21] dmem/dout0[22] dmem/dout0[23] dmem/dout0[24] dmem/dout0[25] dmem/dout0[26]
+ dmem/dout0[27] dmem/dout0[28] dmem/dout0[29] dmem/dout0[30] dmem/dout0[31] la_data_out[0]
+ la_data_out[1] la_data_out[2] la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[30] la_data_out[31] vccd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
.ends

