VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_interface
  CLASS BLOCK ;
  FOREIGN wb_interface ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 152.360 200.000 152.960 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 155.760 200.000 156.360 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 159.160 200.000 159.760 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 162.560 200.000 163.160 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 165.960 200.000 166.560 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 169.360 200.000 169.960 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 172.760 200.000 173.360 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.160 200.000 176.760 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 179.560 200.000 180.160 ;
    END
  END addr0[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 19.760 200.000 20.360 ;
    END
  END clk0
  PIN csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 23.160 200.000 23.760 ;
    END
  END csb0
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 43.560 200.000 44.160 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 77.560 200.000 78.160 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 80.960 200.000 81.560 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 84.360 200.000 84.960 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 87.760 200.000 88.360 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 91.160 200.000 91.760 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 94.560 200.000 95.160 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 97.960 200.000 98.560 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 101.360 200.000 101.960 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 104.760 200.000 105.360 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 108.160 200.000 108.760 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 46.960 200.000 47.560 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 111.560 200.000 112.160 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 114.960 200.000 115.560 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 118.360 200.000 118.960 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 121.760 200.000 122.360 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.160 200.000 125.760 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 128.560 200.000 129.160 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 131.960 200.000 132.560 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 135.360 200.000 135.960 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 138.760 200.000 139.360 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 142.160 200.000 142.760 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 50.360 200.000 50.960 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 145.560 200.000 146.160 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.960 200.000 149.560 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 53.760 200.000 54.360 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 57.160 200.000 57.760 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 60.560 200.000 61.160 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 63.960 200.000 64.560 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 67.360 200.000 67.960 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 70.760 200.000 71.360 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.160 200.000 74.760 ;
    END
  END din0[9]
  PIN imem_rd_cs1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 16.360 200.000 16.960 ;
    END
  END imem_rd_cs1
  PIN processor_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 182.960 200.000 183.560 ;
    END
  END processor_reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END wbs_dat_i[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END wbs_we_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 26.560 200.000 27.160 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 29.960 200.000 30.560 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 33.360 200.000 33.960 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 36.760 200.000 37.360 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 40.160 200.000 40.760 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 187.920 ;
      LAYER met2 ;
        RECT 6.530 10.695 191.720 187.865 ;
      LAYER met3 ;
        RECT 4.000 183.960 196.000 187.845 ;
        RECT 4.000 182.560 195.600 183.960 ;
        RECT 4.000 180.560 196.000 182.560 ;
        RECT 4.000 179.160 195.600 180.560 ;
        RECT 4.000 177.160 196.000 179.160 ;
        RECT 4.000 175.760 195.600 177.160 ;
        RECT 4.000 175.120 196.000 175.760 ;
        RECT 4.400 173.760 196.000 175.120 ;
        RECT 4.400 173.720 195.600 173.760 ;
        RECT 4.000 173.080 195.600 173.720 ;
        RECT 4.400 172.360 195.600 173.080 ;
        RECT 4.400 171.680 196.000 172.360 ;
        RECT 4.000 171.040 196.000 171.680 ;
        RECT 4.400 170.360 196.000 171.040 ;
        RECT 4.400 169.640 195.600 170.360 ;
        RECT 4.000 169.000 195.600 169.640 ;
        RECT 4.400 168.960 195.600 169.000 ;
        RECT 4.400 167.600 196.000 168.960 ;
        RECT 4.000 166.960 196.000 167.600 ;
        RECT 4.400 165.560 195.600 166.960 ;
        RECT 4.000 164.920 196.000 165.560 ;
        RECT 4.400 163.560 196.000 164.920 ;
        RECT 4.400 163.520 195.600 163.560 ;
        RECT 4.000 162.880 195.600 163.520 ;
        RECT 4.400 162.160 195.600 162.880 ;
        RECT 4.400 161.480 196.000 162.160 ;
        RECT 4.000 160.840 196.000 161.480 ;
        RECT 4.400 160.160 196.000 160.840 ;
        RECT 4.400 159.440 195.600 160.160 ;
        RECT 4.000 158.800 195.600 159.440 ;
        RECT 4.400 158.760 195.600 158.800 ;
        RECT 4.400 157.400 196.000 158.760 ;
        RECT 4.000 156.760 196.000 157.400 ;
        RECT 4.400 155.360 195.600 156.760 ;
        RECT 4.000 154.720 196.000 155.360 ;
        RECT 4.400 153.360 196.000 154.720 ;
        RECT 4.400 153.320 195.600 153.360 ;
        RECT 4.000 152.680 195.600 153.320 ;
        RECT 4.400 151.960 195.600 152.680 ;
        RECT 4.400 151.280 196.000 151.960 ;
        RECT 4.000 150.640 196.000 151.280 ;
        RECT 4.400 149.960 196.000 150.640 ;
        RECT 4.400 149.240 195.600 149.960 ;
        RECT 4.000 148.600 195.600 149.240 ;
        RECT 4.400 148.560 195.600 148.600 ;
        RECT 4.400 147.200 196.000 148.560 ;
        RECT 4.000 146.560 196.000 147.200 ;
        RECT 4.400 145.160 195.600 146.560 ;
        RECT 4.000 144.520 196.000 145.160 ;
        RECT 4.400 143.160 196.000 144.520 ;
        RECT 4.400 143.120 195.600 143.160 ;
        RECT 4.000 142.480 195.600 143.120 ;
        RECT 4.400 141.760 195.600 142.480 ;
        RECT 4.400 141.080 196.000 141.760 ;
        RECT 4.000 140.440 196.000 141.080 ;
        RECT 4.400 139.760 196.000 140.440 ;
        RECT 4.400 139.040 195.600 139.760 ;
        RECT 4.000 138.400 195.600 139.040 ;
        RECT 4.400 138.360 195.600 138.400 ;
        RECT 4.400 137.000 196.000 138.360 ;
        RECT 4.000 136.360 196.000 137.000 ;
        RECT 4.400 134.960 195.600 136.360 ;
        RECT 4.000 134.320 196.000 134.960 ;
        RECT 4.400 132.960 196.000 134.320 ;
        RECT 4.400 132.920 195.600 132.960 ;
        RECT 4.000 132.280 195.600 132.920 ;
        RECT 4.400 131.560 195.600 132.280 ;
        RECT 4.400 130.880 196.000 131.560 ;
        RECT 4.000 130.240 196.000 130.880 ;
        RECT 4.400 129.560 196.000 130.240 ;
        RECT 4.400 128.840 195.600 129.560 ;
        RECT 4.000 128.200 195.600 128.840 ;
        RECT 4.400 128.160 195.600 128.200 ;
        RECT 4.400 126.800 196.000 128.160 ;
        RECT 4.000 126.160 196.000 126.800 ;
        RECT 4.400 124.760 195.600 126.160 ;
        RECT 4.000 124.120 196.000 124.760 ;
        RECT 4.400 122.760 196.000 124.120 ;
        RECT 4.400 122.720 195.600 122.760 ;
        RECT 4.000 122.080 195.600 122.720 ;
        RECT 4.400 121.360 195.600 122.080 ;
        RECT 4.400 120.680 196.000 121.360 ;
        RECT 4.000 120.040 196.000 120.680 ;
        RECT 4.400 119.360 196.000 120.040 ;
        RECT 4.400 118.640 195.600 119.360 ;
        RECT 4.000 118.000 195.600 118.640 ;
        RECT 4.400 117.960 195.600 118.000 ;
        RECT 4.400 116.600 196.000 117.960 ;
        RECT 4.000 115.960 196.000 116.600 ;
        RECT 4.400 114.560 195.600 115.960 ;
        RECT 4.000 113.920 196.000 114.560 ;
        RECT 4.400 112.560 196.000 113.920 ;
        RECT 4.400 112.520 195.600 112.560 ;
        RECT 4.000 111.880 195.600 112.520 ;
        RECT 4.400 111.160 195.600 111.880 ;
        RECT 4.400 110.480 196.000 111.160 ;
        RECT 4.000 109.840 196.000 110.480 ;
        RECT 4.400 109.160 196.000 109.840 ;
        RECT 4.400 108.440 195.600 109.160 ;
        RECT 4.000 107.800 195.600 108.440 ;
        RECT 4.400 107.760 195.600 107.800 ;
        RECT 4.400 106.400 196.000 107.760 ;
        RECT 4.000 105.760 196.000 106.400 ;
        RECT 4.400 104.360 195.600 105.760 ;
        RECT 4.000 103.720 196.000 104.360 ;
        RECT 4.400 102.360 196.000 103.720 ;
        RECT 4.400 102.320 195.600 102.360 ;
        RECT 4.000 101.680 195.600 102.320 ;
        RECT 4.400 100.960 195.600 101.680 ;
        RECT 4.400 100.280 196.000 100.960 ;
        RECT 4.000 99.640 196.000 100.280 ;
        RECT 4.400 98.960 196.000 99.640 ;
        RECT 4.400 98.240 195.600 98.960 ;
        RECT 4.000 97.600 195.600 98.240 ;
        RECT 4.400 97.560 195.600 97.600 ;
        RECT 4.400 96.200 196.000 97.560 ;
        RECT 4.000 95.560 196.000 96.200 ;
        RECT 4.400 94.160 195.600 95.560 ;
        RECT 4.000 93.520 196.000 94.160 ;
        RECT 4.400 92.160 196.000 93.520 ;
        RECT 4.400 92.120 195.600 92.160 ;
        RECT 4.000 91.480 195.600 92.120 ;
        RECT 4.400 90.760 195.600 91.480 ;
        RECT 4.400 90.080 196.000 90.760 ;
        RECT 4.000 89.440 196.000 90.080 ;
        RECT 4.400 88.760 196.000 89.440 ;
        RECT 4.400 88.040 195.600 88.760 ;
        RECT 4.000 87.400 195.600 88.040 ;
        RECT 4.400 87.360 195.600 87.400 ;
        RECT 4.400 86.000 196.000 87.360 ;
        RECT 4.000 85.360 196.000 86.000 ;
        RECT 4.400 83.960 195.600 85.360 ;
        RECT 4.000 83.320 196.000 83.960 ;
        RECT 4.400 81.960 196.000 83.320 ;
        RECT 4.400 81.920 195.600 81.960 ;
        RECT 4.000 81.280 195.600 81.920 ;
        RECT 4.400 80.560 195.600 81.280 ;
        RECT 4.400 79.880 196.000 80.560 ;
        RECT 4.000 79.240 196.000 79.880 ;
        RECT 4.400 78.560 196.000 79.240 ;
        RECT 4.400 77.840 195.600 78.560 ;
        RECT 4.000 77.200 195.600 77.840 ;
        RECT 4.400 77.160 195.600 77.200 ;
        RECT 4.400 75.800 196.000 77.160 ;
        RECT 4.000 75.160 196.000 75.800 ;
        RECT 4.400 73.760 195.600 75.160 ;
        RECT 4.000 73.120 196.000 73.760 ;
        RECT 4.400 71.760 196.000 73.120 ;
        RECT 4.400 71.720 195.600 71.760 ;
        RECT 4.000 71.080 195.600 71.720 ;
        RECT 4.400 70.360 195.600 71.080 ;
        RECT 4.400 69.680 196.000 70.360 ;
        RECT 4.000 69.040 196.000 69.680 ;
        RECT 4.400 68.360 196.000 69.040 ;
        RECT 4.400 67.640 195.600 68.360 ;
        RECT 4.000 67.000 195.600 67.640 ;
        RECT 4.400 66.960 195.600 67.000 ;
        RECT 4.400 65.600 196.000 66.960 ;
        RECT 4.000 64.960 196.000 65.600 ;
        RECT 4.400 63.560 195.600 64.960 ;
        RECT 4.000 62.920 196.000 63.560 ;
        RECT 4.400 61.560 196.000 62.920 ;
        RECT 4.400 61.520 195.600 61.560 ;
        RECT 4.000 60.880 195.600 61.520 ;
        RECT 4.400 60.160 195.600 60.880 ;
        RECT 4.400 59.480 196.000 60.160 ;
        RECT 4.000 58.840 196.000 59.480 ;
        RECT 4.400 58.160 196.000 58.840 ;
        RECT 4.400 57.440 195.600 58.160 ;
        RECT 4.000 56.800 195.600 57.440 ;
        RECT 4.400 56.760 195.600 56.800 ;
        RECT 4.400 55.400 196.000 56.760 ;
        RECT 4.000 54.760 196.000 55.400 ;
        RECT 4.400 53.360 195.600 54.760 ;
        RECT 4.000 52.720 196.000 53.360 ;
        RECT 4.400 51.360 196.000 52.720 ;
        RECT 4.400 51.320 195.600 51.360 ;
        RECT 4.000 50.680 195.600 51.320 ;
        RECT 4.400 49.960 195.600 50.680 ;
        RECT 4.400 49.280 196.000 49.960 ;
        RECT 4.000 48.640 196.000 49.280 ;
        RECT 4.400 47.960 196.000 48.640 ;
        RECT 4.400 47.240 195.600 47.960 ;
        RECT 4.000 46.600 195.600 47.240 ;
        RECT 4.400 46.560 195.600 46.600 ;
        RECT 4.400 45.200 196.000 46.560 ;
        RECT 4.000 44.560 196.000 45.200 ;
        RECT 4.400 43.160 195.600 44.560 ;
        RECT 4.000 42.520 196.000 43.160 ;
        RECT 4.400 41.160 196.000 42.520 ;
        RECT 4.400 41.120 195.600 41.160 ;
        RECT 4.000 40.480 195.600 41.120 ;
        RECT 4.400 39.760 195.600 40.480 ;
        RECT 4.400 39.080 196.000 39.760 ;
        RECT 4.000 38.440 196.000 39.080 ;
        RECT 4.400 37.760 196.000 38.440 ;
        RECT 4.400 37.040 195.600 37.760 ;
        RECT 4.000 36.400 195.600 37.040 ;
        RECT 4.400 36.360 195.600 36.400 ;
        RECT 4.400 35.000 196.000 36.360 ;
        RECT 4.000 34.360 196.000 35.000 ;
        RECT 4.400 32.960 195.600 34.360 ;
        RECT 4.000 32.320 196.000 32.960 ;
        RECT 4.400 30.960 196.000 32.320 ;
        RECT 4.400 30.920 195.600 30.960 ;
        RECT 4.000 30.280 195.600 30.920 ;
        RECT 4.400 29.560 195.600 30.280 ;
        RECT 4.400 28.880 196.000 29.560 ;
        RECT 4.000 28.240 196.000 28.880 ;
        RECT 4.400 27.560 196.000 28.240 ;
        RECT 4.400 26.840 195.600 27.560 ;
        RECT 4.000 26.200 195.600 26.840 ;
        RECT 4.400 26.160 195.600 26.200 ;
        RECT 4.400 24.800 196.000 26.160 ;
        RECT 4.000 24.160 196.000 24.800 ;
        RECT 4.000 22.760 195.600 24.160 ;
        RECT 4.000 20.760 196.000 22.760 ;
        RECT 4.000 19.360 195.600 20.760 ;
        RECT 4.000 17.360 196.000 19.360 ;
        RECT 4.000 15.960 195.600 17.360 ;
        RECT 4.000 10.715 196.000 15.960 ;
      LAYER met4 ;
        RECT 13.175 120.535 13.505 138.545 ;
  END
END wb_interface
END LIBRARY

