magic
tech sky130B
magscale 1 2
timestamp 1661333511
<< viali >>
rect 37841 36737 37875 36771
rect 38025 36601 38059 36635
rect 37381 36533 37415 36567
rect 37381 36125 37415 36159
rect 37841 36125 37875 36159
rect 1409 35989 1443 36023
rect 38025 35989 38059 36023
rect 1409 35649 1443 35683
rect 37381 35649 37415 35683
rect 37841 35649 37875 35683
rect 2053 35513 2087 35547
rect 1593 35445 1627 35479
rect 38025 35445 38059 35479
rect 1409 35037 1443 35071
rect 37381 35037 37415 35071
rect 37841 35037 37875 35071
rect 1593 34901 1627 34935
rect 2053 34901 2087 34935
rect 38025 34901 38059 34935
rect 1409 34561 1443 34595
rect 2237 34561 2271 34595
rect 2697 34561 2731 34595
rect 1593 34357 1627 34391
rect 2053 34357 2087 34391
rect 1409 33949 1443 33983
rect 2605 33949 2639 33983
rect 37841 33949 37875 33983
rect 1593 33813 1627 33847
rect 2053 33813 2087 33847
rect 37289 33813 37323 33847
rect 38025 33813 38059 33847
rect 1409 33473 1443 33507
rect 3065 33473 3099 33507
rect 37841 33473 37875 33507
rect 1593 33337 1627 33371
rect 2605 33269 2639 33303
rect 37381 33269 37415 33303
rect 38025 33269 38059 33303
rect 1777 33065 1811 33099
rect 2697 32997 2731 33031
rect 2145 32929 2179 32963
rect 1685 32861 1719 32895
rect 2053 32861 2087 32895
rect 2881 32861 2915 32895
rect 37841 32861 37875 32895
rect 1501 32725 1535 32759
rect 37381 32725 37415 32759
rect 38025 32725 38059 32759
rect 2881 32521 2915 32555
rect 1409 32385 1443 32419
rect 2053 32385 2087 32419
rect 2237 32385 2271 32419
rect 3065 32385 3099 32419
rect 3525 32385 3559 32419
rect 37381 32385 37415 32419
rect 37841 32385 37875 32419
rect 2329 32249 2363 32283
rect 1593 32181 1627 32215
rect 38025 32181 38059 32215
rect 1593 31909 1627 31943
rect 1409 31773 1443 31807
rect 2605 31773 2639 31807
rect 2053 31705 2087 31739
rect 1409 31297 1443 31331
rect 2237 31297 2271 31331
rect 2697 31297 2731 31331
rect 37381 31297 37415 31331
rect 37841 31297 37875 31331
rect 38025 31161 38059 31195
rect 1593 31093 1627 31127
rect 2053 31093 2087 31127
rect 1961 30889 1995 30923
rect 2053 30753 2087 30787
rect 1869 30685 1903 30719
rect 2145 30685 2179 30719
rect 19901 30685 19935 30719
rect 20545 30685 20579 30719
rect 37841 30685 37875 30719
rect 2605 30617 2639 30651
rect 1685 30549 1719 30583
rect 20085 30549 20119 30583
rect 37381 30549 37415 30583
rect 38025 30549 38059 30583
rect 37289 30277 37323 30311
rect 1409 30209 1443 30243
rect 2053 30209 2087 30243
rect 2697 30209 2731 30243
rect 37841 30209 37875 30243
rect 1593 30073 1627 30107
rect 2237 30005 2271 30039
rect 38025 30005 38059 30039
rect 2053 29801 2087 29835
rect 1409 29597 1443 29631
rect 2237 29597 2271 29631
rect 2697 29597 2731 29631
rect 19993 29597 20027 29631
rect 20637 29597 20671 29631
rect 37841 29597 37875 29631
rect 3801 29529 3835 29563
rect 1593 29461 1627 29495
rect 20177 29461 20211 29495
rect 38025 29461 38059 29495
rect 1593 29257 1627 29291
rect 1409 29121 1443 29155
rect 2605 29121 2639 29155
rect 20085 29121 20119 29155
rect 20729 29121 20763 29155
rect 2053 29053 2087 29087
rect 20269 28985 20303 29019
rect 37289 28713 37323 28747
rect 1409 28509 1443 28543
rect 19993 28509 20027 28543
rect 20637 28509 20671 28543
rect 37841 28509 37875 28543
rect 2053 28441 2087 28475
rect 1593 28373 1627 28407
rect 20177 28373 20211 28407
rect 38025 28373 38059 28407
rect 37289 28169 37323 28203
rect 1409 28033 1443 28067
rect 2237 28033 2271 28067
rect 2697 28033 2731 28067
rect 19901 28033 19935 28067
rect 20545 28033 20579 28067
rect 37841 28033 37875 28067
rect 20085 27897 20119 27931
rect 1593 27829 1627 27863
rect 2053 27829 2087 27863
rect 38025 27829 38059 27863
rect 37289 27557 37323 27591
rect 1409 27421 1443 27455
rect 2605 27421 2639 27455
rect 37841 27421 37875 27455
rect 1593 27285 1627 27319
rect 2053 27285 2087 27319
rect 38025 27285 38059 27319
rect 1685 27013 1719 27047
rect 1961 26945 1995 26979
rect 19901 26945 19935 26979
rect 20545 26945 20579 26979
rect 37841 26945 37875 26979
rect 1777 26877 1811 26911
rect 20085 26809 20119 26843
rect 1961 26741 1995 26775
rect 2145 26741 2179 26775
rect 2697 26741 2731 26775
rect 38025 26741 38059 26775
rect 2697 26537 2731 26571
rect 1593 26469 1627 26503
rect 20453 26401 20487 26435
rect 1409 26333 1443 26367
rect 2053 26333 2087 26367
rect 2881 26333 2915 26367
rect 19809 26333 19843 26367
rect 2237 26197 2271 26231
rect 19993 26197 20027 26231
rect 2605 25993 2639 26027
rect 37289 25993 37323 26027
rect 1409 25857 1443 25891
rect 3157 25857 3191 25891
rect 19625 25857 19659 25891
rect 20269 25857 20303 25891
rect 37841 25857 37875 25891
rect 19809 25721 19843 25755
rect 38025 25721 38059 25755
rect 1593 25653 1627 25687
rect 2053 25653 2087 25687
rect 37289 25449 37323 25483
rect 1409 25245 1443 25279
rect 2605 25245 2639 25279
rect 19625 25245 19659 25279
rect 20269 25245 20303 25279
rect 37841 25245 37875 25279
rect 1593 25109 1627 25143
rect 2145 25109 2179 25143
rect 19809 25109 19843 25143
rect 38025 25109 38059 25143
rect 1409 24769 1443 24803
rect 2237 24769 2271 24803
rect 37289 24769 37323 24803
rect 37841 24769 37875 24803
rect 1593 24633 1627 24667
rect 2053 24565 2087 24599
rect 2789 24565 2823 24599
rect 38025 24565 38059 24599
rect 1685 24361 1719 24395
rect 1777 24225 1811 24259
rect 1685 24157 1719 24191
rect 1961 24157 1995 24191
rect 2789 24157 2823 24191
rect 19809 24157 19843 24191
rect 20453 24157 20487 24191
rect 37841 24157 37875 24191
rect 2145 24021 2179 24055
rect 2605 24021 2639 24055
rect 19993 24021 20027 24055
rect 38025 24021 38059 24055
rect 1593 23817 1627 23851
rect 2237 23749 2271 23783
rect 1409 23681 1443 23715
rect 2421 23681 2455 23715
rect 2513 23681 2547 23715
rect 19993 23681 20027 23715
rect 20637 23681 20671 23715
rect 20177 23545 20211 23579
rect 2237 23477 2271 23511
rect 2697 23477 2731 23511
rect 37289 23273 37323 23307
rect 2605 23205 2639 23239
rect 1409 23069 1443 23103
rect 2053 23069 2087 23103
rect 4261 23069 4295 23103
rect 20177 23069 20211 23103
rect 20821 23069 20855 23103
rect 37841 23069 37875 23103
rect 1593 22933 1627 22967
rect 4353 22933 4387 22967
rect 20361 22933 20395 22967
rect 38025 22933 38059 22967
rect 1409 22593 1443 22627
rect 2053 22593 2087 22627
rect 20177 22593 20211 22627
rect 20821 22593 20855 22627
rect 37841 22593 37875 22627
rect 20361 22457 20395 22491
rect 1593 22389 1627 22423
rect 38025 22389 38059 22423
rect 37289 22049 37323 22083
rect 1409 21981 1443 22015
rect 2053 21981 2087 22015
rect 37841 21981 37875 22015
rect 1593 21845 1627 21879
rect 38025 21845 38059 21879
rect 1409 21505 1443 21539
rect 2053 21505 2087 21539
rect 19993 21505 20027 21539
rect 20637 21505 20671 21539
rect 37841 21505 37875 21539
rect 20177 21369 20211 21403
rect 1593 21301 1627 21335
rect 2697 21301 2731 21335
rect 38025 21301 38059 21335
rect 1409 20893 1443 20927
rect 2237 20893 2271 20927
rect 2697 20893 2731 20927
rect 19993 20893 20027 20927
rect 20637 20893 20671 20927
rect 1593 20757 1627 20791
rect 2053 20757 2087 20791
rect 19441 20757 19475 20791
rect 20177 20757 20211 20791
rect 37289 20553 37323 20587
rect 1685 20485 1719 20519
rect 21005 20485 21039 20519
rect 1961 20417 1995 20451
rect 2605 20417 2639 20451
rect 3249 20417 3283 20451
rect 18981 20417 19015 20451
rect 19717 20417 19751 20451
rect 20361 20417 20395 20451
rect 37841 20417 37875 20451
rect 1777 20349 1811 20383
rect 19901 20281 19935 20315
rect 20545 20281 20579 20315
rect 38025 20281 38059 20315
rect 1685 20213 1719 20247
rect 2145 20213 2179 20247
rect 2789 20213 2823 20247
rect 19165 20213 19199 20247
rect 1961 20009 1995 20043
rect 2329 20009 2363 20043
rect 1961 19873 1995 19907
rect 1869 19805 1903 19839
rect 2145 19805 2179 19839
rect 2789 19805 2823 19839
rect 19717 19805 19751 19839
rect 19901 19805 19935 19839
rect 37841 19805 37875 19839
rect 20453 19737 20487 19771
rect 20637 19737 20671 19771
rect 2973 19669 3007 19703
rect 18613 19669 18647 19703
rect 21097 19669 21131 19703
rect 38025 19669 38059 19703
rect 1593 19465 1627 19499
rect 2237 19465 2271 19499
rect 17969 19465 18003 19499
rect 19165 19465 19199 19499
rect 21281 19465 21315 19499
rect 37289 19465 37323 19499
rect 2789 19397 2823 19431
rect 1409 19329 1443 19363
rect 2053 19329 2087 19363
rect 18981 19329 19015 19363
rect 19717 19329 19751 19363
rect 20453 19329 20487 19363
rect 21097 19329 21131 19363
rect 37841 19329 37875 19363
rect 3249 19261 3283 19295
rect 19901 19261 19935 19295
rect 20637 19193 20671 19227
rect 18429 19125 18463 19159
rect 38025 19125 38059 19159
rect 1869 18921 1903 18955
rect 2421 18921 2455 18955
rect 21005 18921 21039 18955
rect 37289 18921 37323 18955
rect 1777 18717 1811 18751
rect 1961 18717 1995 18751
rect 19717 18717 19751 18751
rect 37841 18717 37875 18751
rect 19901 18649 19935 18683
rect 20361 18581 20395 18615
rect 38025 18581 38059 18615
rect 1409 18241 1443 18275
rect 2053 18241 2087 18275
rect 2697 18241 2731 18275
rect 1593 18105 1627 18139
rect 2237 18105 2271 18139
rect 19533 18037 19567 18071
rect 1593 17833 1627 17867
rect 2053 17765 2087 17799
rect 19901 17697 19935 17731
rect 1409 17629 1443 17663
rect 20361 17629 20395 17663
rect 21005 17629 21039 17663
rect 37289 17629 37323 17663
rect 37841 17629 37875 17663
rect 19717 17561 19751 17595
rect 18613 17493 18647 17527
rect 20545 17493 20579 17527
rect 38025 17493 38059 17527
rect 2053 17289 2087 17323
rect 20361 17221 20395 17255
rect 21005 17221 21039 17255
rect 1409 17153 1443 17187
rect 2605 17153 2639 17187
rect 19625 17153 19659 17187
rect 37841 17153 37875 17187
rect 20545 17085 20579 17119
rect 1593 17017 1627 17051
rect 19809 17017 19843 17051
rect 18981 16949 19015 16983
rect 38025 16949 38059 16983
rect 20729 16745 20763 16779
rect 1409 16541 1443 16575
rect 2053 16541 2087 16575
rect 2697 16541 2731 16575
rect 19441 16541 19475 16575
rect 20085 16541 20119 16575
rect 37841 16541 37875 16575
rect 37289 16473 37323 16507
rect 1593 16405 1627 16439
rect 2237 16405 2271 16439
rect 19625 16405 19659 16439
rect 20269 16405 20303 16439
rect 38025 16405 38059 16439
rect 19349 16201 19383 16235
rect 37289 16201 37323 16235
rect 2053 16133 2087 16167
rect 1409 16065 1443 16099
rect 19809 16065 19843 16099
rect 20453 16065 20487 16099
rect 37841 16065 37875 16099
rect 1593 15929 1627 15963
rect 19993 15929 20027 15963
rect 38025 15861 38059 15895
rect 2053 15657 2087 15691
rect 1409 15453 1443 15487
rect 2605 15453 2639 15487
rect 1593 15317 1627 15351
rect 37289 15113 37323 15147
rect 1409 14977 1443 15011
rect 2053 14977 2087 15011
rect 2697 14977 2731 15011
rect 19993 14977 20027 15011
rect 20637 14977 20671 15011
rect 37841 14977 37875 15011
rect 1593 14841 1627 14875
rect 2237 14841 2271 14875
rect 20177 14841 20211 14875
rect 38025 14841 38059 14875
rect 2053 14569 2087 14603
rect 37289 14569 37323 14603
rect 1409 14365 1443 14399
rect 2605 14365 2639 14399
rect 19993 14365 20027 14399
rect 20637 14365 20671 14399
rect 37841 14365 37875 14399
rect 1593 14229 1627 14263
rect 20177 14229 20211 14263
rect 38025 14229 38059 14263
rect 1593 14025 1627 14059
rect 37289 14025 37323 14059
rect 1409 13889 1443 13923
rect 2053 13889 2087 13923
rect 2697 13889 2731 13923
rect 19993 13889 20027 13923
rect 20637 13889 20671 13923
rect 37841 13889 37875 13923
rect 3249 13821 3283 13855
rect 20177 13753 20211 13787
rect 2237 13685 2271 13719
rect 38025 13685 38059 13719
rect 37289 13481 37323 13515
rect 1961 13345 1995 13379
rect 2237 13277 2271 13311
rect 2697 13277 2731 13311
rect 37841 13277 37875 13311
rect 2881 13141 2915 13175
rect 38025 13141 38059 13175
rect 2789 12869 2823 12903
rect 1961 12801 1995 12835
rect 19809 12801 19843 12835
rect 20453 12801 20487 12835
rect 2237 12733 2271 12767
rect 19993 12665 20027 12699
rect 2145 12393 2179 12427
rect 2605 12393 2639 12427
rect 37289 12393 37323 12427
rect 1409 12189 1443 12223
rect 19809 12189 19843 12223
rect 20453 12189 20487 12223
rect 37841 12189 37875 12223
rect 1593 12053 1627 12087
rect 19993 12053 20027 12087
rect 38025 12053 38059 12087
rect 37289 11849 37323 11883
rect 1961 11713 1995 11747
rect 37841 11713 37875 11747
rect 2237 11645 2271 11679
rect 2697 11645 2731 11679
rect 38025 11509 38059 11543
rect 2053 11305 2087 11339
rect 1593 11237 1627 11271
rect 19993 11237 20027 11271
rect 38025 11237 38059 11271
rect 1409 11101 1443 11135
rect 2605 11101 2639 11135
rect 19809 11101 19843 11135
rect 20453 11101 20487 11135
rect 37841 11101 37875 11135
rect 1409 10625 1443 10659
rect 2053 10625 2087 10659
rect 2697 10625 2731 10659
rect 37841 10625 37875 10659
rect 2237 10489 2271 10523
rect 1593 10421 1627 10455
rect 37289 10421 37323 10455
rect 38025 10421 38059 10455
rect 1961 10081 1995 10115
rect 2237 10013 2271 10047
rect 2697 10013 2731 10047
rect 19717 10013 19751 10047
rect 20361 10013 20395 10047
rect 19901 9877 19935 9911
rect 2053 9673 2087 9707
rect 1409 9537 1443 9571
rect 19717 9537 19751 9571
rect 20361 9537 20395 9571
rect 37841 9537 37875 9571
rect 1593 9401 1627 9435
rect 19901 9401 19935 9435
rect 38025 9401 38059 9435
rect 2053 9129 2087 9163
rect 1593 9061 1627 9095
rect 1409 8925 1443 8959
rect 2605 8925 2639 8959
rect 37841 8925 37875 8959
rect 20269 8857 20303 8891
rect 19349 8789 19383 8823
rect 20821 8789 20855 8823
rect 37289 8789 37323 8823
rect 38025 8789 38059 8823
rect 19073 8585 19107 8619
rect 2329 8517 2363 8551
rect 2513 8517 2547 8551
rect 1409 8449 1443 8483
rect 19809 8449 19843 8483
rect 20637 8449 20671 8483
rect 37841 8449 37875 8483
rect 19625 8381 19659 8415
rect 20453 8381 20487 8415
rect 1593 8313 1627 8347
rect 38025 8313 38059 8347
rect 19993 8245 20027 8279
rect 20821 8245 20855 8279
rect 2053 8041 2087 8075
rect 18613 8041 18647 8075
rect 1593 7973 1627 8007
rect 1409 7837 1443 7871
rect 2605 7837 2639 7871
rect 19625 7837 19659 7871
rect 19809 7837 19843 7871
rect 20637 7837 20671 7871
rect 21281 7837 21315 7871
rect 37841 7837 37875 7871
rect 19993 7701 20027 7735
rect 20821 7701 20855 7735
rect 21465 7701 21499 7735
rect 38025 7701 38059 7735
rect 18613 7497 18647 7531
rect 1869 7361 1903 7395
rect 2513 7361 2547 7395
rect 19165 7361 19199 7395
rect 19349 7361 19383 7395
rect 19993 7361 20027 7395
rect 20637 7361 20671 7395
rect 2053 7225 2087 7259
rect 18061 7225 18095 7259
rect 19533 7157 19567 7191
rect 20821 7157 20855 7191
rect 1777 6749 1811 6783
rect 1961 6749 1995 6783
rect 2605 6749 2639 6783
rect 3065 6749 3099 6783
rect 20177 6749 20211 6783
rect 37841 6749 37875 6783
rect 1869 6613 1903 6647
rect 2421 6613 2455 6647
rect 20361 6613 20395 6647
rect 38025 6613 38059 6647
rect 1685 6273 1719 6307
rect 20361 6273 20395 6307
rect 21005 6273 21039 6307
rect 37841 6273 37875 6307
rect 20453 6137 20487 6171
rect 1501 6069 1535 6103
rect 38025 6069 38059 6103
rect 37841 5661 37875 5695
rect 1501 5593 1535 5627
rect 3249 5593 3283 5627
rect 38025 5525 38059 5559
rect 1593 5321 1627 5355
rect 2145 5321 2179 5355
rect 2697 5253 2731 5287
rect 1409 5185 1443 5219
rect 2053 5185 2087 5219
rect 2237 5185 2271 5219
rect 37841 5185 37875 5219
rect 37289 4981 37323 5015
rect 38025 4981 38059 5015
rect 1961 4777 1995 4811
rect 3249 4573 3283 4607
rect 3801 4573 3835 4607
rect 2789 4233 2823 4267
rect 1676 4165 1710 4199
rect 1409 4097 1443 4131
rect 37933 4097 37967 4131
rect 38117 3961 38151 3995
rect 37381 3893 37415 3927
rect 2053 3485 2087 3519
rect 38117 3485 38151 3519
rect 1869 3349 1903 3383
rect 3893 3145 3927 3179
rect 2605 3077 2639 3111
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 37366 36728 37372 36780
rect 37424 36768 37430 36780
rect 37829 36771 37887 36777
rect 37829 36768 37841 36771
rect 37424 36740 37841 36768
rect 37424 36728 37430 36740
rect 37829 36737 37841 36740
rect 37875 36737 37887 36771
rect 37829 36731 37887 36737
rect 38010 36632 38016 36644
rect 37971 36604 38016 36632
rect 38010 36592 38016 36604
rect 38068 36592 38074 36644
rect 37366 36564 37372 36576
rect 37327 36536 37372 36564
rect 37366 36524 37372 36536
rect 37424 36524 37430 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 37369 36159 37427 36165
rect 37369 36125 37381 36159
rect 37415 36156 37427 36159
rect 37829 36159 37887 36165
rect 37829 36156 37841 36159
rect 37415 36128 37841 36156
rect 37415 36125 37427 36128
rect 37369 36119 37427 36125
rect 37829 36125 37841 36128
rect 37875 36156 37887 36159
rect 38194 36156 38200 36168
rect 37875 36128 38200 36156
rect 37875 36125 37887 36128
rect 37829 36119 37887 36125
rect 38194 36116 38200 36128
rect 38252 36116 38258 36168
rect 1394 36020 1400 36032
rect 1355 35992 1400 36020
rect 1394 35980 1400 35992
rect 1452 35980 1458 36032
rect 38010 36020 38016 36032
rect 37971 35992 38016 36020
rect 38010 35980 38016 35992
rect 38068 35980 38074 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1394 35680 1400 35692
rect 1355 35652 1400 35680
rect 1394 35640 1400 35652
rect 1452 35640 1458 35692
rect 37369 35683 37427 35689
rect 37369 35649 37381 35683
rect 37415 35680 37427 35683
rect 37734 35680 37740 35692
rect 37415 35652 37740 35680
rect 37415 35649 37427 35652
rect 37369 35643 37427 35649
rect 37734 35640 37740 35652
rect 37792 35680 37798 35692
rect 37829 35683 37887 35689
rect 37829 35680 37841 35683
rect 37792 35652 37841 35680
rect 37792 35640 37798 35652
rect 37829 35649 37841 35652
rect 37875 35649 37887 35683
rect 37829 35643 37887 35649
rect 1486 35504 1492 35556
rect 1544 35544 1550 35556
rect 2041 35547 2099 35553
rect 2041 35544 2053 35547
rect 1544 35516 2053 35544
rect 1544 35504 1550 35516
rect 2041 35513 2053 35516
rect 2087 35513 2099 35547
rect 2041 35507 2099 35513
rect 1581 35479 1639 35485
rect 1581 35445 1593 35479
rect 1627 35476 1639 35479
rect 2498 35476 2504 35488
rect 1627 35448 2504 35476
rect 1627 35445 1639 35448
rect 1581 35439 1639 35445
rect 2498 35436 2504 35448
rect 2556 35436 2562 35488
rect 38010 35476 38016 35488
rect 37971 35448 38016 35476
rect 38010 35436 38016 35448
rect 38068 35436 38074 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35068 1455 35071
rect 1486 35068 1492 35080
rect 1443 35040 1492 35068
rect 1443 35037 1455 35040
rect 1397 35031 1455 35037
rect 1486 35028 1492 35040
rect 1544 35028 1550 35080
rect 37369 35071 37427 35077
rect 37369 35037 37381 35071
rect 37415 35068 37427 35071
rect 37829 35071 37887 35077
rect 37829 35068 37841 35071
rect 37415 35040 37841 35068
rect 37415 35037 37427 35040
rect 37369 35031 37427 35037
rect 37829 35037 37841 35040
rect 37875 35068 37887 35071
rect 38102 35068 38108 35080
rect 37875 35040 38108 35068
rect 37875 35037 37887 35040
rect 37829 35031 37887 35037
rect 38102 35028 38108 35040
rect 38160 35028 38166 35080
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 2038 34932 2044 34944
rect 1999 34904 2044 34932
rect 2038 34892 2044 34904
rect 2096 34892 2102 34944
rect 38010 34932 38016 34944
rect 37971 34904 38016 34932
rect 38010 34892 38016 34904
rect 38068 34892 38074 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1578 34688 1584 34740
rect 1636 34728 1642 34740
rect 19242 34728 19248 34740
rect 1636 34700 19248 34728
rect 1636 34688 1642 34700
rect 19242 34688 19248 34700
rect 19300 34688 19306 34740
rect 1394 34592 1400 34604
rect 1355 34564 1400 34592
rect 1394 34552 1400 34564
rect 1452 34592 1458 34604
rect 2038 34592 2044 34604
rect 1452 34564 2044 34592
rect 1452 34552 1458 34564
rect 2038 34552 2044 34564
rect 2096 34552 2102 34604
rect 2222 34592 2228 34604
rect 2183 34564 2228 34592
rect 2222 34552 2228 34564
rect 2280 34592 2286 34604
rect 2685 34595 2743 34601
rect 2685 34592 2697 34595
rect 2280 34564 2697 34592
rect 2280 34552 2286 34564
rect 2685 34561 2697 34564
rect 2731 34561 2743 34595
rect 2685 34555 2743 34561
rect 1581 34391 1639 34397
rect 1581 34357 1593 34391
rect 1627 34388 1639 34391
rect 1670 34388 1676 34400
rect 1627 34360 1676 34388
rect 1627 34357 1639 34360
rect 1581 34351 1639 34357
rect 1670 34348 1676 34360
rect 1728 34348 1734 34400
rect 2038 34388 2044 34400
rect 1999 34360 2044 34388
rect 2038 34348 2044 34360
rect 2096 34348 2102 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1394 33980 1400 33992
rect 1355 33952 1400 33980
rect 1394 33940 1400 33952
rect 1452 33980 1458 33992
rect 2593 33983 2651 33989
rect 2593 33980 2605 33983
rect 1452 33952 2605 33980
rect 1452 33940 1458 33952
rect 2593 33949 2605 33952
rect 2639 33949 2651 33983
rect 37829 33983 37887 33989
rect 37829 33980 37841 33983
rect 2593 33943 2651 33949
rect 37292 33952 37841 33980
rect 37292 33856 37320 33952
rect 37829 33949 37841 33952
rect 37875 33949 37887 33983
rect 37829 33943 37887 33949
rect 1578 33844 1584 33856
rect 1539 33816 1584 33844
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 1762 33804 1768 33856
rect 1820 33844 1826 33856
rect 2041 33847 2099 33853
rect 2041 33844 2053 33847
rect 1820 33816 2053 33844
rect 1820 33804 1826 33816
rect 2041 33813 2053 33816
rect 2087 33813 2099 33847
rect 37274 33844 37280 33856
rect 37235 33816 37280 33844
rect 2041 33807 2099 33813
rect 37274 33804 37280 33816
rect 37332 33804 37338 33856
rect 38010 33844 38016 33856
rect 37971 33816 38016 33844
rect 38010 33804 38016 33816
rect 38068 33804 38074 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1578 33600 1584 33652
rect 1636 33640 1642 33652
rect 19150 33640 19156 33652
rect 1636 33612 19156 33640
rect 1636 33600 1642 33612
rect 19150 33600 19156 33612
rect 19208 33600 19214 33652
rect 1397 33507 1455 33513
rect 1397 33473 1409 33507
rect 1443 33504 1455 33507
rect 1578 33504 1584 33516
rect 1443 33476 1584 33504
rect 1443 33473 1455 33476
rect 1397 33467 1455 33473
rect 1578 33464 1584 33476
rect 1636 33504 1642 33516
rect 3053 33507 3111 33513
rect 3053 33504 3065 33507
rect 1636 33476 3065 33504
rect 1636 33464 1642 33476
rect 3053 33473 3065 33476
rect 3099 33473 3111 33507
rect 3053 33467 3111 33473
rect 37458 33464 37464 33516
rect 37516 33504 37522 33516
rect 37829 33507 37887 33513
rect 37829 33504 37841 33507
rect 37516 33476 37841 33504
rect 37516 33464 37522 33476
rect 37829 33473 37841 33476
rect 37875 33473 37887 33507
rect 37829 33467 37887 33473
rect 1581 33371 1639 33377
rect 1581 33337 1593 33371
rect 1627 33368 1639 33371
rect 19978 33368 19984 33380
rect 1627 33340 19984 33368
rect 1627 33337 1639 33340
rect 1581 33331 1639 33337
rect 19978 33328 19984 33340
rect 20036 33328 20042 33380
rect 2593 33303 2651 33309
rect 2593 33269 2605 33303
rect 2639 33300 2651 33303
rect 2866 33300 2872 33312
rect 2639 33272 2872 33300
rect 2639 33269 2651 33272
rect 2593 33263 2651 33269
rect 2866 33260 2872 33272
rect 2924 33260 2930 33312
rect 37369 33303 37427 33309
rect 37369 33269 37381 33303
rect 37415 33300 37427 33303
rect 37458 33300 37464 33312
rect 37415 33272 37464 33300
rect 37415 33269 37427 33272
rect 37369 33263 37427 33269
rect 37458 33260 37464 33272
rect 37516 33260 37522 33312
rect 38010 33300 38016 33312
rect 37971 33272 38016 33300
rect 38010 33260 38016 33272
rect 38068 33260 38074 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1765 33099 1823 33105
rect 1765 33065 1777 33099
rect 1811 33096 1823 33099
rect 2038 33096 2044 33108
rect 1811 33068 2044 33096
rect 1811 33065 1823 33068
rect 1765 33059 1823 33065
rect 2038 33056 2044 33068
rect 2096 33056 2102 33108
rect 2685 33031 2743 33037
rect 2685 33028 2697 33031
rect 2148 33000 2697 33028
rect 2148 32969 2176 33000
rect 2685 32997 2697 33000
rect 2731 32997 2743 33031
rect 2685 32991 2743 32997
rect 2133 32963 2191 32969
rect 2133 32929 2145 32963
rect 2179 32929 2191 32963
rect 2133 32923 2191 32929
rect 1670 32892 1676 32904
rect 1631 32864 1676 32892
rect 1670 32852 1676 32864
rect 1728 32852 1734 32904
rect 2038 32892 2044 32904
rect 1999 32864 2044 32892
rect 2038 32852 2044 32864
rect 2096 32852 2102 32904
rect 2866 32892 2872 32904
rect 2827 32864 2872 32892
rect 2866 32852 2872 32864
rect 2924 32852 2930 32904
rect 37829 32895 37887 32901
rect 37829 32892 37841 32895
rect 37568 32864 37841 32892
rect 37568 32768 37596 32864
rect 37829 32861 37841 32864
rect 37875 32861 37887 32895
rect 37829 32855 37887 32861
rect 1486 32756 1492 32768
rect 1447 32728 1492 32756
rect 1486 32716 1492 32728
rect 1544 32716 1550 32768
rect 37369 32759 37427 32765
rect 37369 32725 37381 32759
rect 37415 32756 37427 32759
rect 37550 32756 37556 32768
rect 37415 32728 37556 32756
rect 37415 32725 37427 32728
rect 37369 32719 37427 32725
rect 37550 32716 37556 32728
rect 37608 32716 37614 32768
rect 38010 32756 38016 32768
rect 37971 32728 38016 32756
rect 38010 32716 38016 32728
rect 38068 32716 38074 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 2038 32512 2044 32564
rect 2096 32552 2102 32564
rect 2869 32555 2927 32561
rect 2869 32552 2881 32555
rect 2096 32524 2881 32552
rect 2096 32512 2102 32524
rect 2869 32521 2881 32524
rect 2915 32521 2927 32555
rect 2869 32515 2927 32521
rect 1762 32484 1768 32496
rect 1412 32456 1768 32484
rect 1412 32425 1440 32456
rect 1762 32444 1768 32456
rect 1820 32444 1826 32496
rect 1397 32419 1455 32425
rect 1397 32385 1409 32419
rect 1443 32385 1455 32419
rect 1397 32379 1455 32385
rect 1486 32376 1492 32428
rect 1544 32416 1550 32428
rect 2041 32419 2099 32425
rect 2041 32416 2053 32419
rect 1544 32388 2053 32416
rect 1544 32376 1550 32388
rect 2041 32385 2053 32388
rect 2087 32416 2099 32419
rect 2130 32416 2136 32428
rect 2087 32388 2136 32416
rect 2087 32385 2099 32388
rect 2041 32379 2099 32385
rect 2130 32376 2136 32388
rect 2188 32376 2194 32428
rect 2225 32419 2283 32425
rect 2225 32385 2237 32419
rect 2271 32385 2283 32419
rect 3050 32416 3056 32428
rect 3011 32388 3056 32416
rect 2225 32379 2283 32385
rect 1854 32308 1860 32360
rect 1912 32348 1918 32360
rect 2240 32348 2268 32379
rect 3050 32376 3056 32388
rect 3108 32416 3114 32428
rect 3513 32419 3571 32425
rect 3513 32416 3525 32419
rect 3108 32388 3525 32416
rect 3108 32376 3114 32388
rect 3513 32385 3525 32388
rect 3559 32385 3571 32419
rect 3513 32379 3571 32385
rect 37369 32419 37427 32425
rect 37369 32385 37381 32419
rect 37415 32416 37427 32419
rect 37829 32419 37887 32425
rect 37829 32416 37841 32419
rect 37415 32388 37841 32416
rect 37415 32385 37427 32388
rect 37369 32379 37427 32385
rect 37829 32385 37841 32388
rect 37875 32416 37887 32419
rect 38286 32416 38292 32428
rect 37875 32388 38292 32416
rect 37875 32385 37887 32388
rect 37829 32379 37887 32385
rect 38286 32376 38292 32388
rect 38344 32376 38350 32428
rect 1912 32320 2268 32348
rect 1912 32308 1918 32320
rect 2317 32283 2375 32289
rect 2317 32249 2329 32283
rect 2363 32280 2375 32283
rect 37366 32280 37372 32292
rect 2363 32252 37372 32280
rect 2363 32249 2375 32252
rect 2317 32243 2375 32249
rect 37366 32240 37372 32252
rect 37424 32240 37430 32292
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 1670 32212 1676 32224
rect 1627 32184 1676 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 1670 32172 1676 32184
rect 1728 32172 1734 32224
rect 38010 32212 38016 32224
rect 37971 32184 38016 32212
rect 38010 32172 38016 32184
rect 38068 32172 38074 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1581 31943 1639 31949
rect 1581 31909 1593 31943
rect 1627 31940 1639 31943
rect 2682 31940 2688 31952
rect 1627 31912 2688 31940
rect 1627 31909 1639 31912
rect 1581 31903 1639 31909
rect 2682 31900 2688 31912
rect 2740 31900 2746 31952
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31804 1458 31816
rect 2593 31807 2651 31813
rect 2593 31804 2605 31807
rect 1452 31776 2605 31804
rect 1452 31764 1458 31776
rect 2593 31773 2605 31776
rect 2639 31773 2651 31807
rect 2593 31767 2651 31773
rect 1486 31696 1492 31748
rect 1544 31736 1550 31748
rect 2041 31739 2099 31745
rect 2041 31736 2053 31739
rect 1544 31708 2053 31736
rect 1544 31696 1550 31708
rect 2041 31705 2053 31708
rect 2087 31705 2099 31739
rect 2041 31699 2099 31705
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1397 31331 1455 31337
rect 1397 31297 1409 31331
rect 1443 31328 1455 31331
rect 1486 31328 1492 31340
rect 1443 31300 1492 31328
rect 1443 31297 1455 31300
rect 1397 31291 1455 31297
rect 1486 31288 1492 31300
rect 1544 31288 1550 31340
rect 2222 31328 2228 31340
rect 2183 31300 2228 31328
rect 2222 31288 2228 31300
rect 2280 31328 2286 31340
rect 2685 31331 2743 31337
rect 2685 31328 2697 31331
rect 2280 31300 2697 31328
rect 2280 31288 2286 31300
rect 2685 31297 2697 31300
rect 2731 31297 2743 31331
rect 2685 31291 2743 31297
rect 37369 31331 37427 31337
rect 37369 31297 37381 31331
rect 37415 31328 37427 31331
rect 37829 31331 37887 31337
rect 37829 31328 37841 31331
rect 37415 31300 37841 31328
rect 37415 31297 37427 31300
rect 37369 31291 37427 31297
rect 37829 31297 37841 31300
rect 37875 31328 37887 31331
rect 37918 31328 37924 31340
rect 37875 31300 37924 31328
rect 37875 31297 37887 31300
rect 37829 31291 37887 31297
rect 37918 31288 37924 31300
rect 37976 31288 37982 31340
rect 38010 31192 38016 31204
rect 37971 31164 38016 31192
rect 38010 31152 38016 31164
rect 38068 31152 38074 31204
rect 1581 31127 1639 31133
rect 1581 31093 1593 31127
rect 1627 31124 1639 31127
rect 1854 31124 1860 31136
rect 1627 31096 1860 31124
rect 1627 31093 1639 31096
rect 1581 31087 1639 31093
rect 1854 31084 1860 31096
rect 1912 31084 1918 31136
rect 2038 31124 2044 31136
rect 1999 31096 2044 31124
rect 2038 31084 2044 31096
rect 2096 31084 2102 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1946 30920 1952 30932
rect 1907 30892 1952 30920
rect 1946 30880 1952 30892
rect 2004 30880 2010 30932
rect 2038 30784 2044 30796
rect 1999 30756 2044 30784
rect 2038 30744 2044 30756
rect 2096 30744 2102 30796
rect 1854 30716 1860 30728
rect 1815 30688 1860 30716
rect 1854 30676 1860 30688
rect 1912 30676 1918 30728
rect 2130 30716 2136 30728
rect 2091 30688 2136 30716
rect 2130 30676 2136 30688
rect 2188 30676 2194 30728
rect 2498 30676 2504 30728
rect 2556 30716 2562 30728
rect 19889 30719 19947 30725
rect 19889 30716 19901 30719
rect 2556 30688 19901 30716
rect 2556 30676 2562 30688
rect 19889 30685 19901 30688
rect 19935 30716 19947 30719
rect 20533 30719 20591 30725
rect 20533 30716 20545 30719
rect 19935 30688 20545 30716
rect 19935 30685 19947 30688
rect 19889 30679 19947 30685
rect 20533 30685 20545 30688
rect 20579 30685 20591 30719
rect 37829 30719 37887 30725
rect 37829 30716 37841 30719
rect 20533 30679 20591 30685
rect 37660 30688 37841 30716
rect 1578 30608 1584 30660
rect 1636 30648 1642 30660
rect 2593 30651 2651 30657
rect 2593 30648 2605 30651
rect 1636 30620 2605 30648
rect 1636 30608 1642 30620
rect 2593 30617 2605 30620
rect 2639 30617 2651 30651
rect 34514 30648 34520 30660
rect 2593 30611 2651 30617
rect 20088 30620 34520 30648
rect 1673 30583 1731 30589
rect 1673 30549 1685 30583
rect 1719 30580 1731 30583
rect 2130 30580 2136 30592
rect 1719 30552 2136 30580
rect 1719 30549 1731 30552
rect 1673 30543 1731 30549
rect 2130 30540 2136 30552
rect 2188 30540 2194 30592
rect 20088 30589 20116 30620
rect 34514 30608 34520 30620
rect 34572 30608 34578 30660
rect 37660 30592 37688 30688
rect 37829 30685 37841 30688
rect 37875 30685 37887 30719
rect 37829 30679 37887 30685
rect 20073 30583 20131 30589
rect 20073 30549 20085 30583
rect 20119 30549 20131 30583
rect 20073 30543 20131 30549
rect 37369 30583 37427 30589
rect 37369 30549 37381 30583
rect 37415 30580 37427 30583
rect 37642 30580 37648 30592
rect 37415 30552 37648 30580
rect 37415 30549 37427 30552
rect 37369 30543 37427 30549
rect 37642 30540 37648 30552
rect 37700 30540 37706 30592
rect 38010 30580 38016 30592
rect 37971 30552 38016 30580
rect 38010 30540 38016 30552
rect 38068 30540 38074 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 34514 30268 34520 30320
rect 34572 30308 34578 30320
rect 37277 30311 37335 30317
rect 37277 30308 37289 30311
rect 34572 30280 37289 30308
rect 34572 30268 34578 30280
rect 37277 30277 37289 30280
rect 37323 30308 37335 30311
rect 37323 30280 37872 30308
rect 37323 30277 37335 30280
rect 37277 30271 37335 30277
rect 1397 30243 1455 30249
rect 1397 30209 1409 30243
rect 1443 30240 1455 30243
rect 1486 30240 1492 30252
rect 1443 30212 1492 30240
rect 1443 30209 1455 30212
rect 1397 30203 1455 30209
rect 1486 30200 1492 30212
rect 1544 30200 1550 30252
rect 2038 30240 2044 30252
rect 1999 30212 2044 30240
rect 2038 30200 2044 30212
rect 2096 30240 2102 30252
rect 37844 30249 37872 30280
rect 2685 30243 2743 30249
rect 2685 30240 2697 30243
rect 2096 30212 2697 30240
rect 2096 30200 2102 30212
rect 2685 30209 2697 30212
rect 2731 30209 2743 30243
rect 2685 30203 2743 30209
rect 37829 30243 37887 30249
rect 37829 30209 37841 30243
rect 37875 30209 37887 30243
rect 37829 30203 37887 30209
rect 1581 30107 1639 30113
rect 1581 30073 1593 30107
rect 1627 30104 1639 30107
rect 2406 30104 2412 30116
rect 1627 30076 2412 30104
rect 1627 30073 1639 30076
rect 1581 30067 1639 30073
rect 2406 30064 2412 30076
rect 2464 30064 2470 30116
rect 2222 30036 2228 30048
rect 2183 30008 2228 30036
rect 2222 29996 2228 30008
rect 2280 29996 2286 30048
rect 38010 30036 38016 30048
rect 37971 30008 38016 30036
rect 38010 29996 38016 30008
rect 38068 29996 38074 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1946 29792 1952 29844
rect 2004 29832 2010 29844
rect 2041 29835 2099 29841
rect 2041 29832 2053 29835
rect 2004 29804 2053 29832
rect 2004 29792 2010 29804
rect 2041 29801 2053 29804
rect 2087 29801 2099 29835
rect 2041 29795 2099 29801
rect 2222 29792 2228 29844
rect 2280 29832 2286 29844
rect 12434 29832 12440 29844
rect 2280 29804 12440 29832
rect 2280 29792 2286 29804
rect 12434 29792 12440 29804
rect 12492 29792 12498 29844
rect 1397 29631 1455 29637
rect 1397 29597 1409 29631
rect 1443 29597 1455 29631
rect 2222 29628 2228 29640
rect 2183 29600 2228 29628
rect 1397 29591 1455 29597
rect 1302 29520 1308 29572
rect 1360 29560 1366 29572
rect 1412 29560 1440 29591
rect 2222 29588 2228 29600
rect 2280 29628 2286 29640
rect 2685 29631 2743 29637
rect 2685 29628 2697 29631
rect 2280 29600 2697 29628
rect 2280 29588 2286 29600
rect 2685 29597 2697 29600
rect 2731 29597 2743 29631
rect 2685 29591 2743 29597
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 19981 29631 20039 29637
rect 19981 29628 19993 29631
rect 19300 29600 19993 29628
rect 19300 29588 19306 29600
rect 19981 29597 19993 29600
rect 20027 29628 20039 29631
rect 20625 29631 20683 29637
rect 20625 29628 20637 29631
rect 20027 29600 20637 29628
rect 20027 29597 20039 29600
rect 19981 29591 20039 29597
rect 20625 29597 20637 29600
rect 20671 29597 20683 29631
rect 37829 29631 37887 29637
rect 37829 29628 37841 29631
rect 20625 29591 20683 29597
rect 26206 29600 37841 29628
rect 3789 29563 3847 29569
rect 3789 29560 3801 29563
rect 1360 29532 3801 29560
rect 1360 29520 1366 29532
rect 3789 29529 3801 29532
rect 3835 29529 3847 29563
rect 26206 29560 26234 29600
rect 37829 29597 37841 29600
rect 37875 29597 37887 29631
rect 37829 29591 37887 29597
rect 3789 29523 3847 29529
rect 20180 29532 26234 29560
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 1762 29492 1768 29504
rect 1627 29464 1768 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 1762 29452 1768 29464
rect 1820 29452 1826 29504
rect 20180 29501 20208 29532
rect 20165 29495 20223 29501
rect 20165 29461 20177 29495
rect 20211 29461 20223 29495
rect 38010 29492 38016 29504
rect 37971 29464 38016 29492
rect 20165 29455 20223 29461
rect 38010 29452 38016 29464
rect 38068 29452 38074 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1581 29291 1639 29297
rect 1581 29257 1593 29291
rect 1627 29288 1639 29291
rect 2498 29288 2504 29300
rect 1627 29260 2504 29288
rect 1627 29257 1639 29260
rect 1581 29251 1639 29257
rect 2498 29248 2504 29260
rect 2556 29248 2562 29300
rect 1394 29152 1400 29164
rect 1355 29124 1400 29152
rect 1394 29112 1400 29124
rect 1452 29152 1458 29164
rect 2593 29155 2651 29161
rect 2593 29152 2605 29155
rect 1452 29124 2605 29152
rect 1452 29112 1458 29124
rect 2593 29121 2605 29124
rect 2639 29121 2651 29155
rect 2593 29115 2651 29121
rect 19150 29112 19156 29164
rect 19208 29152 19214 29164
rect 20073 29155 20131 29161
rect 20073 29152 20085 29155
rect 19208 29124 20085 29152
rect 19208 29112 19214 29124
rect 20073 29121 20085 29124
rect 20119 29152 20131 29155
rect 20717 29155 20775 29161
rect 20717 29152 20729 29155
rect 20119 29124 20729 29152
rect 20119 29121 20131 29124
rect 20073 29115 20131 29121
rect 20717 29121 20729 29124
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 1578 29044 1584 29096
rect 1636 29084 1642 29096
rect 2041 29087 2099 29093
rect 2041 29084 2053 29087
rect 1636 29056 2053 29084
rect 1636 29044 1642 29056
rect 2041 29053 2053 29056
rect 2087 29053 2099 29087
rect 2041 29047 2099 29053
rect 20257 29019 20315 29025
rect 20257 28985 20269 29019
rect 20303 29016 20315 29019
rect 37274 29016 37280 29028
rect 20303 28988 37280 29016
rect 20303 28985 20315 28988
rect 20257 28979 20315 28985
rect 37274 28976 37280 28988
rect 37332 28976 37338 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 37274 28744 37280 28756
rect 37235 28716 37280 28744
rect 37274 28704 37280 28716
rect 37332 28704 37338 28756
rect 1397 28543 1455 28549
rect 1397 28509 1409 28543
rect 1443 28540 1455 28543
rect 1578 28540 1584 28552
rect 1443 28512 1584 28540
rect 1443 28509 1455 28512
rect 1397 28503 1455 28509
rect 1578 28500 1584 28512
rect 1636 28500 1642 28552
rect 19978 28540 19984 28552
rect 19939 28512 19984 28540
rect 19978 28500 19984 28512
rect 20036 28540 20042 28552
rect 20625 28543 20683 28549
rect 20625 28540 20637 28543
rect 20036 28512 20637 28540
rect 20036 28500 20042 28512
rect 20625 28509 20637 28512
rect 20671 28509 20683 28543
rect 20625 28503 20683 28509
rect 37274 28500 37280 28552
rect 37332 28540 37338 28552
rect 37829 28543 37887 28549
rect 37829 28540 37841 28543
rect 37332 28512 37841 28540
rect 37332 28500 37338 28512
rect 37829 28509 37841 28512
rect 37875 28509 37887 28543
rect 37829 28503 37887 28509
rect 1486 28432 1492 28484
rect 1544 28472 1550 28484
rect 2041 28475 2099 28481
rect 2041 28472 2053 28475
rect 1544 28444 2053 28472
rect 1544 28432 1550 28444
rect 2041 28441 2053 28444
rect 2087 28441 2099 28475
rect 37182 28472 37188 28484
rect 2041 28435 2099 28441
rect 20180 28444 37188 28472
rect 1581 28407 1639 28413
rect 1581 28373 1593 28407
rect 1627 28404 1639 28407
rect 2590 28404 2596 28416
rect 1627 28376 2596 28404
rect 1627 28373 1639 28376
rect 1581 28367 1639 28373
rect 2590 28364 2596 28376
rect 2648 28364 2654 28416
rect 20180 28413 20208 28444
rect 37182 28432 37188 28444
rect 37240 28432 37246 28484
rect 20165 28407 20223 28413
rect 20165 28373 20177 28407
rect 20211 28373 20223 28407
rect 38010 28404 38016 28416
rect 37971 28376 38016 28404
rect 20165 28367 20223 28373
rect 38010 28364 38016 28376
rect 38068 28364 38074 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 37182 28160 37188 28212
rect 37240 28200 37246 28212
rect 37277 28203 37335 28209
rect 37277 28200 37289 28203
rect 37240 28172 37289 28200
rect 37240 28160 37246 28172
rect 37277 28169 37289 28172
rect 37323 28169 37335 28203
rect 37277 28163 37335 28169
rect 1670 28092 1676 28144
rect 1728 28132 1734 28144
rect 1728 28104 19932 28132
rect 1728 28092 1734 28104
rect 1397 28067 1455 28073
rect 1397 28033 1409 28067
rect 1443 28064 1455 28067
rect 1486 28064 1492 28076
rect 1443 28036 1492 28064
rect 1443 28033 1455 28036
rect 1397 28027 1455 28033
rect 1486 28024 1492 28036
rect 1544 28024 1550 28076
rect 2222 28064 2228 28076
rect 2183 28036 2228 28064
rect 2222 28024 2228 28036
rect 2280 28064 2286 28076
rect 19904 28073 19932 28104
rect 2685 28067 2743 28073
rect 2685 28064 2697 28067
rect 2280 28036 2697 28064
rect 2280 28024 2286 28036
rect 2685 28033 2697 28036
rect 2731 28033 2743 28067
rect 2685 28027 2743 28033
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28064 19947 28067
rect 20533 28067 20591 28073
rect 20533 28064 20545 28067
rect 19935 28036 20545 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 20533 28033 20545 28036
rect 20579 28033 20591 28067
rect 37292 28064 37320 28163
rect 37829 28067 37887 28073
rect 37829 28064 37841 28067
rect 37292 28036 37841 28064
rect 20533 28027 20591 28033
rect 37829 28033 37841 28036
rect 37875 28033 37887 28067
rect 37829 28027 37887 28033
rect 37274 27996 37280 28008
rect 26206 27968 37280 27996
rect 20073 27931 20131 27937
rect 20073 27897 20085 27931
rect 20119 27928 20131 27931
rect 26206 27928 26234 27968
rect 37274 27956 37280 27968
rect 37332 27956 37338 28008
rect 20119 27900 26234 27928
rect 20119 27897 20131 27900
rect 20073 27891 20131 27897
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 1946 27860 1952 27872
rect 1627 27832 1952 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 1946 27820 1952 27832
rect 2004 27820 2010 27872
rect 2038 27820 2044 27872
rect 2096 27860 2102 27872
rect 38010 27860 38016 27872
rect 2096 27832 2141 27860
rect 37971 27832 38016 27860
rect 2096 27820 2102 27832
rect 38010 27820 38016 27832
rect 38068 27820 38074 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 37274 27588 37280 27600
rect 37235 27560 37280 27588
rect 37274 27548 37280 27560
rect 37332 27548 37338 27600
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27452 1458 27464
rect 2593 27455 2651 27461
rect 2593 27452 2605 27455
rect 1452 27424 2605 27452
rect 1452 27412 1458 27424
rect 2593 27421 2605 27424
rect 2639 27421 2651 27455
rect 37292 27452 37320 27548
rect 37829 27455 37887 27461
rect 37829 27452 37841 27455
rect 37292 27424 37841 27452
rect 2593 27415 2651 27421
rect 37829 27421 37841 27424
rect 37875 27421 37887 27455
rect 37829 27415 37887 27421
rect 1596 27356 6914 27384
rect 1596 27325 1624 27356
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27285 1639 27319
rect 1581 27279 1639 27285
rect 1670 27276 1676 27328
rect 1728 27316 1734 27328
rect 2041 27319 2099 27325
rect 2041 27316 2053 27319
rect 1728 27288 2053 27316
rect 1728 27276 1734 27288
rect 2041 27285 2053 27288
rect 2087 27285 2099 27319
rect 6886 27316 6914 27356
rect 19426 27316 19432 27328
rect 6886 27288 19432 27316
rect 2041 27279 2099 27285
rect 19426 27276 19432 27288
rect 19484 27276 19490 27328
rect 38010 27316 38016 27328
rect 37971 27288 38016 27316
rect 38010 27276 38016 27288
rect 38068 27276 38074 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1673 27047 1731 27053
rect 1673 27013 1685 27047
rect 1719 27044 1731 27047
rect 2038 27044 2044 27056
rect 1719 27016 2044 27044
rect 1719 27013 1731 27016
rect 1673 27007 1731 27013
rect 2038 27004 2044 27016
rect 2096 27004 2102 27056
rect 1946 26976 1952 26988
rect 1907 26948 1952 26976
rect 1946 26936 1952 26948
rect 2004 26936 2010 26988
rect 19889 26979 19947 26985
rect 19889 26976 19901 26979
rect 6886 26948 19901 26976
rect 1762 26908 1768 26920
rect 1723 26880 1768 26908
rect 1762 26868 1768 26880
rect 1820 26868 1826 26920
rect 2682 26868 2688 26920
rect 2740 26908 2746 26920
rect 6886 26908 6914 26948
rect 19889 26945 19901 26948
rect 19935 26976 19947 26979
rect 20533 26979 20591 26985
rect 20533 26976 20545 26979
rect 19935 26948 20545 26976
rect 19935 26945 19947 26948
rect 19889 26939 19947 26945
rect 20533 26945 20545 26948
rect 20579 26945 20591 26979
rect 37829 26979 37887 26985
rect 37829 26976 37841 26979
rect 20533 26939 20591 26945
rect 26206 26948 37841 26976
rect 2740 26880 6914 26908
rect 2740 26868 2746 26880
rect 20073 26843 20131 26849
rect 20073 26809 20085 26843
rect 20119 26840 20131 26843
rect 26206 26840 26234 26948
rect 37829 26945 37841 26948
rect 37875 26945 37887 26979
rect 37829 26939 37887 26945
rect 20119 26812 26234 26840
rect 20119 26809 20131 26812
rect 20073 26803 20131 26809
rect 1946 26772 1952 26784
rect 1907 26744 1952 26772
rect 1946 26732 1952 26744
rect 2004 26732 2010 26784
rect 2130 26772 2136 26784
rect 2091 26744 2136 26772
rect 2130 26732 2136 26744
rect 2188 26732 2194 26784
rect 2685 26775 2743 26781
rect 2685 26741 2697 26775
rect 2731 26772 2743 26775
rect 2774 26772 2780 26784
rect 2731 26744 2780 26772
rect 2731 26741 2743 26744
rect 2685 26735 2743 26741
rect 2774 26732 2780 26744
rect 2832 26732 2838 26784
rect 38010 26772 38016 26784
rect 37971 26744 38016 26772
rect 38010 26732 38016 26744
rect 38068 26732 38074 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1946 26528 1952 26580
rect 2004 26568 2010 26580
rect 2685 26571 2743 26577
rect 2685 26568 2697 26571
rect 2004 26540 2697 26568
rect 2004 26528 2010 26540
rect 2685 26537 2697 26540
rect 2731 26537 2743 26571
rect 2685 26531 2743 26537
rect 1581 26503 1639 26509
rect 1581 26469 1593 26503
rect 1627 26500 1639 26503
rect 1762 26500 1768 26512
rect 1627 26472 1768 26500
rect 1627 26469 1639 26472
rect 1581 26463 1639 26469
rect 1762 26460 1768 26472
rect 1820 26460 1826 26512
rect 2590 26392 2596 26444
rect 2648 26432 2654 26444
rect 20441 26435 20499 26441
rect 20441 26432 20453 26435
rect 2648 26404 2912 26432
rect 2648 26392 2654 26404
rect 1397 26367 1455 26373
rect 1397 26333 1409 26367
rect 1443 26364 1455 26367
rect 1486 26364 1492 26376
rect 1443 26336 1492 26364
rect 1443 26333 1455 26336
rect 1397 26327 1455 26333
rect 1486 26324 1492 26336
rect 1544 26364 1550 26376
rect 1670 26364 1676 26376
rect 1544 26336 1676 26364
rect 1544 26324 1550 26336
rect 1670 26324 1676 26336
rect 1728 26324 1734 26376
rect 2038 26364 2044 26376
rect 1951 26336 2044 26364
rect 2038 26324 2044 26336
rect 2096 26364 2102 26376
rect 2774 26364 2780 26376
rect 2096 26336 2780 26364
rect 2096 26324 2102 26336
rect 2774 26324 2780 26336
rect 2832 26324 2838 26376
rect 2884 26373 2912 26404
rect 19812 26404 20453 26432
rect 2869 26367 2927 26373
rect 2869 26333 2881 26367
rect 2915 26333 2927 26367
rect 2869 26327 2927 26333
rect 12434 26324 12440 26376
rect 12492 26364 12498 26376
rect 19812 26373 19840 26404
rect 20441 26401 20453 26404
rect 20487 26401 20499 26435
rect 20441 26395 20499 26401
rect 19797 26367 19855 26373
rect 19797 26364 19809 26367
rect 12492 26336 19809 26364
rect 12492 26324 12498 26336
rect 19797 26333 19809 26336
rect 19843 26333 19855 26367
rect 19797 26327 19855 26333
rect 19996 26336 26234 26364
rect 16574 26296 16580 26308
rect 2240 26268 16580 26296
rect 2240 26237 2268 26268
rect 16574 26256 16580 26268
rect 16632 26256 16638 26308
rect 19996 26237 20024 26336
rect 26206 26296 26234 26336
rect 37182 26296 37188 26308
rect 26206 26268 37188 26296
rect 37182 26256 37188 26268
rect 37240 26256 37246 26308
rect 2225 26231 2283 26237
rect 2225 26197 2237 26231
rect 2271 26228 2283 26231
rect 19981 26231 20039 26237
rect 2271 26200 2305 26228
rect 2271 26197 2283 26200
rect 2225 26191 2283 26197
rect 19981 26197 19993 26231
rect 20027 26228 20039 26231
rect 20027 26200 20061 26228
rect 20027 26197 20039 26200
rect 19981 26191 20039 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 2590 26024 2596 26036
rect 2551 25996 2596 26024
rect 2590 25984 2596 25996
rect 2648 25984 2654 26036
rect 37182 25984 37188 26036
rect 37240 26024 37246 26036
rect 37277 26027 37335 26033
rect 37277 26024 37289 26027
rect 37240 25996 37289 26024
rect 37240 25984 37246 25996
rect 37277 25993 37289 25996
rect 37323 25993 37335 26027
rect 37277 25987 37335 25993
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25888 1458 25900
rect 3145 25891 3203 25897
rect 3145 25888 3157 25891
rect 1452 25860 3157 25888
rect 1452 25848 1458 25860
rect 3145 25857 3157 25860
rect 3191 25857 3203 25891
rect 19613 25891 19671 25897
rect 19613 25888 19625 25891
rect 3145 25851 3203 25857
rect 6886 25860 19625 25888
rect 2406 25712 2412 25764
rect 2464 25752 2470 25764
rect 6886 25752 6914 25860
rect 19613 25857 19625 25860
rect 19659 25888 19671 25891
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 19659 25860 20269 25888
rect 19659 25857 19671 25860
rect 19613 25851 19671 25857
rect 20257 25857 20269 25860
rect 20303 25857 20315 25891
rect 37292 25888 37320 25987
rect 37829 25891 37887 25897
rect 37829 25888 37841 25891
rect 37292 25860 37841 25888
rect 20257 25851 20315 25857
rect 37829 25857 37841 25860
rect 37875 25857 37887 25891
rect 37829 25851 37887 25857
rect 2464 25724 6914 25752
rect 19797 25755 19855 25761
rect 2464 25712 2470 25724
rect 19797 25721 19809 25755
rect 19843 25752 19855 25755
rect 37182 25752 37188 25764
rect 19843 25724 37188 25752
rect 19843 25721 19855 25724
rect 19797 25715 19855 25721
rect 37182 25712 37188 25724
rect 37240 25712 37246 25764
rect 38010 25752 38016 25764
rect 37971 25724 38016 25752
rect 38010 25712 38016 25724
rect 38068 25712 38074 25764
rect 1578 25684 1584 25696
rect 1539 25656 1584 25684
rect 1578 25644 1584 25656
rect 1636 25644 1642 25696
rect 1946 25644 1952 25696
rect 2004 25684 2010 25696
rect 2041 25687 2099 25693
rect 2041 25684 2053 25687
rect 2004 25656 2053 25684
rect 2004 25644 2010 25656
rect 2041 25653 2053 25656
rect 2087 25653 2099 25687
rect 2041 25647 2099 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 1578 25440 1584 25492
rect 1636 25480 1642 25492
rect 13814 25480 13820 25492
rect 1636 25452 13820 25480
rect 1636 25440 1642 25452
rect 13814 25440 13820 25452
rect 13872 25440 13878 25492
rect 37182 25440 37188 25492
rect 37240 25480 37246 25492
rect 37277 25483 37335 25489
rect 37277 25480 37289 25483
rect 37240 25452 37289 25480
rect 37240 25440 37246 25452
rect 37277 25449 37289 25452
rect 37323 25449 37335 25483
rect 37277 25443 37335 25449
rect 1397 25279 1455 25285
rect 1397 25245 1409 25279
rect 1443 25276 1455 25279
rect 1486 25276 1492 25288
rect 1443 25248 1492 25276
rect 1443 25245 1455 25248
rect 1397 25239 1455 25245
rect 1486 25236 1492 25248
rect 1544 25276 1550 25288
rect 2593 25279 2651 25285
rect 2593 25276 2605 25279
rect 1544 25248 2605 25276
rect 1544 25236 1550 25248
rect 2593 25245 2605 25248
rect 2639 25245 2651 25279
rect 2593 25239 2651 25245
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25276 19671 25279
rect 20257 25279 20315 25285
rect 20257 25276 20269 25279
rect 19659 25248 20269 25276
rect 19659 25245 19671 25248
rect 19613 25239 19671 25245
rect 20257 25245 20269 25248
rect 20303 25245 20315 25279
rect 37292 25276 37320 25443
rect 37829 25279 37887 25285
rect 37829 25276 37841 25279
rect 37292 25248 37841 25276
rect 20257 25239 20315 25245
rect 37829 25245 37841 25248
rect 37875 25245 37887 25279
rect 37829 25239 37887 25245
rect 2498 25168 2504 25220
rect 2556 25208 2562 25220
rect 19628 25208 19656 25239
rect 33134 25208 33140 25220
rect 2556 25180 19656 25208
rect 19812 25180 33140 25208
rect 2556 25168 2562 25180
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 2130 25140 2136 25152
rect 2091 25112 2136 25140
rect 2130 25100 2136 25112
rect 2188 25100 2194 25152
rect 19812 25149 19840 25180
rect 33134 25168 33140 25180
rect 33192 25168 33198 25220
rect 19797 25143 19855 25149
rect 19797 25109 19809 25143
rect 19843 25109 19855 25143
rect 38010 25140 38016 25152
rect 37971 25112 38016 25140
rect 19797 25103 19855 25109
rect 38010 25100 38016 25112
rect 38068 25100 38074 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1578 24896 1584 24948
rect 1636 24936 1642 24948
rect 19978 24936 19984 24948
rect 1636 24908 19984 24936
rect 1636 24896 1642 24908
rect 19978 24896 19984 24908
rect 20036 24896 20042 24948
rect 1394 24800 1400 24812
rect 1355 24772 1400 24800
rect 1394 24760 1400 24772
rect 1452 24800 1458 24812
rect 1946 24800 1952 24812
rect 1452 24772 1952 24800
rect 1452 24760 1458 24772
rect 1946 24760 1952 24772
rect 2004 24760 2010 24812
rect 2130 24760 2136 24812
rect 2188 24800 2194 24812
rect 2225 24803 2283 24809
rect 2225 24800 2237 24803
rect 2188 24772 2237 24800
rect 2188 24760 2194 24772
rect 2225 24769 2237 24772
rect 2271 24769 2283 24803
rect 2225 24763 2283 24769
rect 33134 24760 33140 24812
rect 33192 24800 33198 24812
rect 37277 24803 37335 24809
rect 37277 24800 37289 24803
rect 33192 24772 37289 24800
rect 33192 24760 33198 24772
rect 37277 24769 37289 24772
rect 37323 24800 37335 24803
rect 37829 24803 37887 24809
rect 37829 24800 37841 24803
rect 37323 24772 37841 24800
rect 37323 24769 37335 24772
rect 37277 24763 37335 24769
rect 37829 24769 37841 24772
rect 37875 24769 37887 24803
rect 37829 24763 37887 24769
rect 1581 24667 1639 24673
rect 1581 24633 1593 24667
rect 1627 24664 1639 24667
rect 1627 24636 6914 24664
rect 1627 24633 1639 24636
rect 1581 24627 1639 24633
rect 1670 24556 1676 24608
rect 1728 24596 1734 24608
rect 2041 24599 2099 24605
rect 2041 24596 2053 24599
rect 1728 24568 2053 24596
rect 1728 24556 1734 24568
rect 2041 24565 2053 24568
rect 2087 24565 2099 24599
rect 2774 24596 2780 24608
rect 2735 24568 2780 24596
rect 2041 24559 2099 24565
rect 2774 24556 2780 24568
rect 2832 24556 2838 24608
rect 6886 24596 6914 24636
rect 17770 24596 17776 24608
rect 6886 24568 17776 24596
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 38010 24596 38016 24608
rect 37971 24568 38016 24596
rect 38010 24556 38016 24568
rect 38068 24556 38074 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1578 24352 1584 24404
rect 1636 24392 1642 24404
rect 1673 24395 1731 24401
rect 1673 24392 1685 24395
rect 1636 24364 1685 24392
rect 1636 24352 1642 24364
rect 1673 24361 1685 24364
rect 1719 24361 1731 24395
rect 1673 24355 1731 24361
rect 1762 24256 1768 24268
rect 1723 24228 1768 24256
rect 1762 24216 1768 24228
rect 1820 24216 1826 24268
rect 1670 24188 1676 24200
rect 1631 24160 1676 24188
rect 1670 24148 1676 24160
rect 1728 24148 1734 24200
rect 1949 24191 2007 24197
rect 1949 24157 1961 24191
rect 1995 24188 2007 24191
rect 2774 24188 2780 24200
rect 1995 24160 2636 24188
rect 2735 24160 2780 24188
rect 1995 24157 2007 24160
rect 1949 24151 2007 24157
rect 2133 24055 2191 24061
rect 2133 24021 2145 24055
rect 2179 24052 2191 24055
rect 2406 24052 2412 24064
rect 2179 24024 2412 24052
rect 2179 24021 2191 24024
rect 2133 24015 2191 24021
rect 2406 24012 2412 24024
rect 2464 24012 2470 24064
rect 2608 24061 2636 24160
rect 2774 24148 2780 24160
rect 2832 24148 2838 24200
rect 19794 24188 19800 24200
rect 19755 24160 19800 24188
rect 19794 24148 19800 24160
rect 19852 24188 19858 24200
rect 20441 24191 20499 24197
rect 20441 24188 20453 24191
rect 19852 24160 20453 24188
rect 19852 24148 19858 24160
rect 20441 24157 20453 24160
rect 20487 24157 20499 24191
rect 37829 24191 37887 24197
rect 37829 24188 37841 24191
rect 20441 24151 20499 24157
rect 26206 24160 37841 24188
rect 26206 24120 26234 24160
rect 37829 24157 37841 24160
rect 37875 24157 37887 24191
rect 37829 24151 37887 24157
rect 19996 24092 26234 24120
rect 19996 24061 20024 24092
rect 2593 24055 2651 24061
rect 2593 24021 2605 24055
rect 2639 24021 2651 24055
rect 2593 24015 2651 24021
rect 19981 24055 20039 24061
rect 19981 24021 19993 24055
rect 20027 24021 20039 24055
rect 38010 24052 38016 24064
rect 37971 24024 38016 24052
rect 19981 24015 20039 24021
rect 38010 24012 38016 24024
rect 38068 24012 38074 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 2222 23780 2228 23792
rect 2183 23752 2228 23780
rect 2222 23740 2228 23752
rect 2280 23740 2286 23792
rect 1397 23715 1455 23721
rect 1397 23681 1409 23715
rect 1443 23712 1455 23715
rect 1486 23712 1492 23724
rect 1443 23684 1492 23712
rect 1443 23681 1455 23684
rect 1397 23675 1455 23681
rect 1486 23672 1492 23684
rect 1544 23672 1550 23724
rect 2406 23712 2412 23724
rect 2367 23684 2412 23712
rect 2406 23672 2412 23684
rect 2464 23672 2470 23724
rect 2498 23672 2504 23724
rect 2556 23712 2562 23724
rect 2556 23684 2601 23712
rect 2556 23672 2562 23684
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 19981 23715 20039 23721
rect 19981 23712 19993 23715
rect 19484 23684 19993 23712
rect 19484 23672 19490 23684
rect 19981 23681 19993 23684
rect 20027 23712 20039 23715
rect 20625 23715 20683 23721
rect 20625 23712 20637 23715
rect 20027 23684 20637 23712
rect 20027 23681 20039 23684
rect 19981 23675 20039 23681
rect 20625 23681 20637 23684
rect 20671 23681 20683 23715
rect 20625 23675 20683 23681
rect 20165 23579 20223 23585
rect 20165 23545 20177 23579
rect 20211 23576 20223 23579
rect 20211 23548 26234 23576
rect 20211 23545 20223 23548
rect 20165 23539 20223 23545
rect 2038 23468 2044 23520
rect 2096 23508 2102 23520
rect 2225 23511 2283 23517
rect 2225 23508 2237 23511
rect 2096 23480 2237 23508
rect 2096 23468 2102 23480
rect 2225 23477 2237 23480
rect 2271 23477 2283 23511
rect 2225 23471 2283 23477
rect 2685 23511 2743 23517
rect 2685 23477 2697 23511
rect 2731 23508 2743 23511
rect 4614 23508 4620 23520
rect 2731 23480 4620 23508
rect 2731 23477 2743 23480
rect 2685 23471 2743 23477
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 26206 23508 26234 23548
rect 37274 23508 37280 23520
rect 26206 23480 37280 23508
rect 37274 23468 37280 23480
rect 37332 23468 37338 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 37274 23304 37280 23316
rect 37235 23276 37280 23304
rect 37274 23264 37280 23276
rect 37332 23264 37338 23316
rect 1486 23196 1492 23248
rect 1544 23236 1550 23248
rect 2593 23239 2651 23245
rect 2593 23236 2605 23239
rect 1544 23208 2605 23236
rect 1544 23196 1550 23208
rect 2593 23205 2605 23208
rect 2639 23205 2651 23239
rect 2593 23199 2651 23205
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23100 1458 23112
rect 2041 23103 2099 23109
rect 2041 23100 2053 23103
rect 1452 23072 2053 23100
rect 1452 23060 1458 23072
rect 2041 23069 2053 23072
rect 2087 23069 2099 23103
rect 2041 23063 2099 23069
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4614 23100 4620 23112
rect 4295 23072 4620 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 16574 23060 16580 23112
rect 16632 23100 16638 23112
rect 20165 23103 20223 23109
rect 20165 23100 20177 23103
rect 16632 23072 20177 23100
rect 16632 23060 16638 23072
rect 20165 23069 20177 23072
rect 20211 23100 20223 23103
rect 20809 23103 20867 23109
rect 20809 23100 20821 23103
rect 20211 23072 20821 23100
rect 20211 23069 20223 23072
rect 20165 23063 20223 23069
rect 20809 23069 20821 23072
rect 20855 23069 20867 23103
rect 20809 23063 20867 23069
rect 37274 23060 37280 23112
rect 37332 23100 37338 23112
rect 37829 23103 37887 23109
rect 37829 23100 37841 23103
rect 37332 23072 37841 23100
rect 37332 23060 37338 23072
rect 37829 23069 37841 23072
rect 37875 23069 37887 23103
rect 37829 23063 37887 23069
rect 31018 23032 31024 23044
rect 20364 23004 31024 23032
rect 1578 22964 1584 22976
rect 1539 22936 1584 22964
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 4341 22967 4399 22973
rect 4341 22933 4353 22967
rect 4387 22964 4399 22967
rect 4614 22964 4620 22976
rect 4387 22936 4620 22964
rect 4387 22933 4399 22936
rect 4341 22927 4399 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 20364 22973 20392 23004
rect 31018 22992 31024 23004
rect 31076 22992 31082 23044
rect 20349 22967 20407 22973
rect 20349 22933 20361 22967
rect 20395 22933 20407 22967
rect 38010 22964 38016 22976
rect 37971 22936 38016 22964
rect 20349 22927 20407 22933
rect 38010 22924 38016 22936
rect 38068 22924 38074 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1578 22720 1584 22772
rect 1636 22760 1642 22772
rect 17862 22760 17868 22772
rect 1636 22732 17868 22760
rect 1636 22720 1642 22732
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22624 1458 22636
rect 2041 22627 2099 22633
rect 2041 22624 2053 22627
rect 1452 22596 2053 22624
rect 1452 22584 1458 22596
rect 2041 22593 2053 22596
rect 2087 22593 2099 22627
rect 2041 22587 2099 22593
rect 13814 22584 13820 22636
rect 13872 22624 13878 22636
rect 20165 22627 20223 22633
rect 20165 22624 20177 22627
rect 13872 22596 20177 22624
rect 13872 22584 13878 22596
rect 20165 22593 20177 22596
rect 20211 22624 20223 22627
rect 20809 22627 20867 22633
rect 20809 22624 20821 22627
rect 20211 22596 20821 22624
rect 20211 22593 20223 22596
rect 20165 22587 20223 22593
rect 20809 22593 20821 22596
rect 20855 22593 20867 22627
rect 20809 22587 20867 22593
rect 31018 22584 31024 22636
rect 31076 22624 31082 22636
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 31076 22596 37841 22624
rect 31076 22584 31082 22596
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 20349 22491 20407 22497
rect 20349 22457 20361 22491
rect 20395 22488 20407 22491
rect 20395 22460 26234 22488
rect 20395 22457 20407 22460
rect 20349 22451 20407 22457
rect 1581 22423 1639 22429
rect 1581 22389 1593 22423
rect 1627 22420 1639 22423
rect 1762 22420 1768 22432
rect 1627 22392 1768 22420
rect 1627 22389 1639 22392
rect 1581 22383 1639 22389
rect 1762 22380 1768 22392
rect 1820 22380 1826 22432
rect 26206 22420 26234 22460
rect 37274 22420 37280 22432
rect 26206 22392 37280 22420
rect 37274 22380 37280 22392
rect 37332 22380 37338 22432
rect 38010 22420 38016 22432
rect 37971 22392 38016 22420
rect 38010 22380 38016 22392
rect 38068 22380 38074 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 37274 22080 37280 22092
rect 37235 22052 37280 22080
rect 37274 22040 37280 22052
rect 37332 22080 37338 22092
rect 37332 22052 37872 22080
rect 37332 22040 37338 22052
rect 1394 22012 1400 22024
rect 1355 21984 1400 22012
rect 1394 21972 1400 21984
rect 1452 22012 1458 22024
rect 37844 22021 37872 22052
rect 2041 22015 2099 22021
rect 2041 22012 2053 22015
rect 1452 21984 2053 22012
rect 1452 21972 1458 21984
rect 2041 21981 2053 21984
rect 2087 21981 2099 22015
rect 2041 21975 2099 21981
rect 37829 22015 37887 22021
rect 37829 21981 37841 22015
rect 37875 21981 37887 22015
rect 37829 21975 37887 21981
rect 1596 21916 6914 21944
rect 1596 21885 1624 21916
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21845 1639 21879
rect 6886 21876 6914 21916
rect 17954 21876 17960 21888
rect 6886 21848 17960 21876
rect 1581 21839 1639 21845
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 38010 21876 38016 21888
rect 37971 21848 38016 21876
rect 38010 21836 38016 21848
rect 38068 21836 38074 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21536 1458 21548
rect 2041 21539 2099 21545
rect 2041 21536 2053 21539
rect 1452 21508 2053 21536
rect 1452 21496 1458 21508
rect 2041 21505 2053 21508
rect 2087 21505 2099 21539
rect 19978 21536 19984 21548
rect 19939 21508 19984 21536
rect 2041 21499 2099 21505
rect 19978 21496 19984 21508
rect 20036 21536 20042 21548
rect 20625 21539 20683 21545
rect 20625 21536 20637 21539
rect 20036 21508 20637 21536
rect 20036 21496 20042 21508
rect 20625 21505 20637 21508
rect 20671 21505 20683 21539
rect 37829 21539 37887 21545
rect 37829 21536 37841 21539
rect 20625 21499 20683 21505
rect 26206 21508 37841 21536
rect 20165 21403 20223 21409
rect 20165 21369 20177 21403
rect 20211 21400 20223 21403
rect 26206 21400 26234 21508
rect 37829 21505 37841 21508
rect 37875 21505 37887 21539
rect 37829 21499 37887 21505
rect 20211 21372 26234 21400
rect 20211 21369 20223 21372
rect 20165 21363 20223 21369
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 2685 21335 2743 21341
rect 2685 21301 2697 21335
rect 2731 21332 2743 21335
rect 2774 21332 2780 21344
rect 2731 21304 2780 21332
rect 2731 21301 2743 21304
rect 2685 21295 2743 21301
rect 2774 21292 2780 21304
rect 2832 21292 2838 21344
rect 38010 21332 38016 21344
rect 37971 21304 38016 21332
rect 38010 21292 38016 21304
rect 38068 21292 38074 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1486 20952 1492 21004
rect 1544 20992 1550 21004
rect 2774 20992 2780 21004
rect 1544 20964 2780 20992
rect 1544 20952 1550 20964
rect 2774 20952 2780 20964
rect 2832 20952 2838 21004
rect 1397 20927 1455 20933
rect 1397 20893 1409 20927
rect 1443 20924 1455 20927
rect 1504 20924 1532 20952
rect 2222 20924 2228 20936
rect 1443 20896 1532 20924
rect 2183 20896 2228 20924
rect 1443 20893 1455 20896
rect 1397 20887 1455 20893
rect 2222 20884 2228 20896
rect 2280 20924 2286 20936
rect 2685 20927 2743 20933
rect 2685 20924 2697 20927
rect 2280 20896 2697 20924
rect 2280 20884 2286 20896
rect 2685 20893 2697 20896
rect 2731 20893 2743 20927
rect 2685 20887 2743 20893
rect 17770 20884 17776 20936
rect 17828 20924 17834 20936
rect 19981 20927 20039 20933
rect 19981 20924 19993 20927
rect 17828 20896 19993 20924
rect 17828 20884 17834 20896
rect 19981 20893 19993 20896
rect 20027 20924 20039 20927
rect 20625 20927 20683 20933
rect 20625 20924 20637 20927
rect 20027 20896 20637 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 20625 20893 20637 20896
rect 20671 20893 20683 20927
rect 20625 20887 20683 20893
rect 18966 20856 18972 20868
rect 1596 20828 18972 20856
rect 1596 20797 1624 20828
rect 18966 20816 18972 20828
rect 19024 20816 19030 20868
rect 33134 20856 33140 20868
rect 20180 20828 33140 20856
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20757 1639 20791
rect 1581 20751 1639 20757
rect 1946 20748 1952 20800
rect 2004 20788 2010 20800
rect 2041 20791 2099 20797
rect 2041 20788 2053 20791
rect 2004 20760 2053 20788
rect 2004 20748 2010 20760
rect 2041 20757 2053 20760
rect 2087 20757 2099 20791
rect 19426 20788 19432 20800
rect 19387 20760 19432 20788
rect 2041 20751 2099 20757
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 20180 20797 20208 20828
rect 33134 20816 33140 20828
rect 33192 20816 33198 20868
rect 20165 20791 20223 20797
rect 20165 20757 20177 20791
rect 20211 20757 20223 20791
rect 20165 20751 20223 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 33134 20544 33140 20596
rect 33192 20584 33198 20596
rect 37277 20587 37335 20593
rect 37277 20584 37289 20587
rect 33192 20556 37289 20584
rect 33192 20544 33198 20556
rect 37277 20553 37289 20556
rect 37323 20553 37335 20587
rect 37277 20547 37335 20553
rect 1578 20476 1584 20528
rect 1636 20516 1642 20528
rect 1673 20519 1731 20525
rect 1673 20516 1685 20519
rect 1636 20488 1685 20516
rect 1636 20476 1642 20488
rect 1673 20485 1685 20488
rect 1719 20485 1731 20519
rect 1673 20479 1731 20485
rect 17862 20476 17868 20528
rect 17920 20516 17926 20528
rect 20993 20519 21051 20525
rect 20993 20516 21005 20519
rect 17920 20488 21005 20516
rect 17920 20476 17926 20488
rect 1946 20448 1952 20460
rect 1907 20420 1952 20448
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 2593 20451 2651 20457
rect 2593 20417 2605 20451
rect 2639 20448 2651 20451
rect 2866 20448 2872 20460
rect 2639 20420 2872 20448
rect 2639 20417 2651 20420
rect 2593 20411 2651 20417
rect 2866 20408 2872 20420
rect 2924 20448 2930 20460
rect 3237 20451 3295 20457
rect 3237 20448 3249 20451
rect 2924 20420 3249 20448
rect 2924 20408 2930 20420
rect 3237 20417 3249 20420
rect 3283 20417 3295 20451
rect 18966 20448 18972 20460
rect 18927 20420 18972 20448
rect 3237 20411 3295 20417
rect 18966 20408 18972 20420
rect 19024 20408 19030 20460
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 20364 20457 20392 20488
rect 20993 20485 21005 20488
rect 21039 20485 21051 20519
rect 20993 20479 21051 20485
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 19484 20420 19717 20448
rect 19484 20408 19490 20420
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 37292 20448 37320 20547
rect 37829 20451 37887 20457
rect 37829 20448 37841 20451
rect 37292 20420 37841 20448
rect 20349 20411 20407 20417
rect 37829 20417 37841 20420
rect 37875 20417 37887 20451
rect 37829 20411 37887 20417
rect 1762 20380 1768 20392
rect 1723 20352 1768 20380
rect 1762 20340 1768 20352
rect 1820 20340 1826 20392
rect 19886 20312 19892 20324
rect 19847 20284 19892 20312
rect 19886 20272 19892 20284
rect 19944 20272 19950 20324
rect 20533 20315 20591 20321
rect 20533 20281 20545 20315
rect 20579 20312 20591 20315
rect 31018 20312 31024 20324
rect 20579 20284 31024 20312
rect 20579 20281 20591 20284
rect 20533 20275 20591 20281
rect 31018 20272 31024 20284
rect 31076 20272 31082 20324
rect 38010 20312 38016 20324
rect 37971 20284 38016 20312
rect 38010 20272 38016 20284
rect 38068 20272 38074 20324
rect 1578 20204 1584 20256
rect 1636 20244 1642 20256
rect 1673 20247 1731 20253
rect 1673 20244 1685 20247
rect 1636 20216 1685 20244
rect 1636 20204 1642 20216
rect 1673 20213 1685 20216
rect 1719 20213 1731 20247
rect 1673 20207 1731 20213
rect 2038 20204 2044 20256
rect 2096 20244 2102 20256
rect 2133 20247 2191 20253
rect 2133 20244 2145 20247
rect 2096 20216 2145 20244
rect 2096 20204 2102 20216
rect 2133 20213 2145 20216
rect 2179 20213 2191 20247
rect 2774 20244 2780 20256
rect 2735 20216 2780 20244
rect 2133 20207 2191 20213
rect 2774 20204 2780 20216
rect 2832 20204 2838 20256
rect 19150 20244 19156 20256
rect 19111 20216 19156 20244
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 2317 20043 2375 20049
rect 2317 20009 2329 20043
rect 2363 20040 2375 20043
rect 2498 20040 2504 20052
rect 2363 20012 2504 20040
rect 2363 20009 2375 20012
rect 2317 20003 2375 20009
rect 2498 20000 2504 20012
rect 2556 20000 2562 20052
rect 19150 20000 19156 20052
rect 19208 20040 19214 20052
rect 31754 20040 31760 20052
rect 19208 20012 31760 20040
rect 19208 20000 19214 20012
rect 31754 20000 31760 20012
rect 31812 20000 31818 20052
rect 2774 19932 2780 19984
rect 2832 19972 2838 19984
rect 21082 19972 21088 19984
rect 2832 19944 21088 19972
rect 2832 19932 2838 19944
rect 21082 19932 21088 19944
rect 21140 19932 21146 19984
rect 1762 19864 1768 19916
rect 1820 19904 1826 19916
rect 1949 19907 2007 19913
rect 1949 19904 1961 19907
rect 1820 19876 1961 19904
rect 1820 19864 1826 19876
rect 1949 19873 1961 19876
rect 1995 19873 2007 19907
rect 1949 19867 2007 19873
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19836 1915 19839
rect 2038 19836 2044 19848
rect 1903 19808 2044 19836
rect 1903 19805 1915 19808
rect 1857 19799 1915 19805
rect 2038 19796 2044 19808
rect 2096 19796 2102 19848
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19836 2191 19839
rect 2222 19836 2228 19848
rect 2179 19808 2228 19836
rect 2179 19805 2191 19808
rect 2133 19799 2191 19805
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 2774 19836 2780 19848
rect 2735 19808 2780 19836
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 18506 19796 18512 19848
rect 18564 19836 18570 19848
rect 19705 19839 19763 19845
rect 19705 19836 19717 19839
rect 18564 19808 19717 19836
rect 18564 19796 18570 19808
rect 19705 19805 19717 19808
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 19935 19808 26234 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 14458 19728 14464 19780
rect 14516 19768 14522 19780
rect 20441 19771 20499 19777
rect 14516 19740 19656 19768
rect 14516 19728 14522 19740
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19700 3019 19703
rect 17862 19700 17868 19712
rect 3007 19672 17868 19700
rect 3007 19669 3019 19672
rect 2961 19663 3019 19669
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 18506 19660 18512 19712
rect 18564 19700 18570 19712
rect 18601 19703 18659 19709
rect 18601 19700 18613 19703
rect 18564 19672 18613 19700
rect 18564 19660 18570 19672
rect 18601 19669 18613 19672
rect 18647 19669 18659 19703
rect 19628 19700 19656 19740
rect 20441 19737 20453 19771
rect 20487 19737 20499 19771
rect 20622 19768 20628 19780
rect 20583 19740 20628 19768
rect 20441 19731 20499 19737
rect 20456 19700 20484 19731
rect 20622 19728 20628 19740
rect 20680 19728 20686 19780
rect 21085 19703 21143 19709
rect 21085 19700 21097 19703
rect 19628 19672 21097 19700
rect 18601 19663 18659 19669
rect 21085 19669 21097 19672
rect 21131 19669 21143 19703
rect 26206 19700 26234 19808
rect 31018 19796 31024 19848
rect 31076 19836 31082 19848
rect 37829 19839 37887 19845
rect 37829 19836 37841 19839
rect 31076 19808 37841 19836
rect 31076 19796 31082 19808
rect 37829 19805 37841 19808
rect 37875 19805 37887 19839
rect 37829 19799 37887 19805
rect 37642 19700 37648 19712
rect 26206 19672 37648 19700
rect 21085 19663 21143 19669
rect 37642 19660 37648 19672
rect 37700 19660 37706 19712
rect 38010 19700 38016 19712
rect 37971 19672 38016 19700
rect 38010 19660 38016 19672
rect 38068 19660 38074 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 2222 19496 2228 19508
rect 2183 19468 2228 19496
rect 2222 19456 2228 19468
rect 2280 19456 2286 19508
rect 17954 19496 17960 19508
rect 17915 19468 17960 19496
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 19153 19499 19211 19505
rect 19153 19465 19165 19499
rect 19199 19465 19211 19499
rect 19153 19459 19211 19465
rect 21269 19499 21327 19505
rect 21269 19465 21281 19499
rect 21315 19496 21327 19499
rect 27522 19496 27528 19508
rect 21315 19468 27528 19496
rect 21315 19465 21327 19468
rect 21269 19459 21327 19465
rect 2774 19428 2780 19440
rect 1412 19400 2360 19428
rect 2735 19400 2780 19428
rect 1412 19372 1440 19400
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 2038 19360 2044 19372
rect 1999 19332 2044 19360
rect 2038 19320 2044 19332
rect 2096 19320 2102 19372
rect 2332 19360 2360 19400
rect 2774 19388 2780 19400
rect 2832 19388 2838 19440
rect 17972 19360 18000 19456
rect 19168 19428 19196 19459
rect 27522 19456 27528 19468
rect 27580 19456 27586 19508
rect 37277 19499 37335 19505
rect 37277 19496 37289 19499
rect 35866 19468 37289 19496
rect 35866 19428 35894 19468
rect 37277 19465 37289 19468
rect 37323 19465 37335 19499
rect 37277 19459 37335 19465
rect 19168 19400 35894 19428
rect 18969 19363 19027 19369
rect 18969 19360 18981 19363
rect 2332 19332 3280 19360
rect 17972 19332 18981 19360
rect 3252 19301 3280 19332
rect 18969 19329 18981 19332
rect 19015 19329 19027 19363
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 18969 19323 19027 19329
rect 19076 19332 19717 19360
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19261 3295 19295
rect 19076 19292 19104 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 20346 19320 20352 19372
rect 20404 19360 20410 19372
rect 20441 19363 20499 19369
rect 20441 19360 20453 19363
rect 20404 19332 20453 19360
rect 20404 19320 20410 19332
rect 20441 19329 20453 19332
rect 20487 19329 20499 19363
rect 21082 19360 21088 19372
rect 21043 19332 21088 19360
rect 20441 19323 20499 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 37292 19360 37320 19459
rect 37829 19363 37887 19369
rect 37829 19360 37841 19363
rect 37292 19332 37841 19360
rect 37829 19329 37841 19332
rect 37875 19329 37887 19363
rect 37829 19323 37887 19329
rect 3237 19255 3295 19261
rect 18432 19264 19104 19292
rect 19889 19295 19947 19301
rect 18432 19168 18460 19264
rect 19889 19261 19901 19295
rect 19935 19292 19947 19295
rect 19935 19264 26234 19292
rect 19935 19261 19947 19264
rect 19889 19255 19947 19261
rect 20625 19227 20683 19233
rect 20625 19193 20637 19227
rect 20671 19224 20683 19227
rect 26206 19224 26234 19264
rect 38286 19224 38292 19236
rect 20671 19196 23428 19224
rect 26206 19196 38292 19224
rect 20671 19193 20683 19196
rect 20625 19187 20683 19193
rect 18414 19156 18420 19168
rect 18375 19128 18420 19156
rect 18414 19116 18420 19128
rect 18472 19116 18478 19168
rect 23400 19156 23428 19196
rect 38286 19184 38292 19196
rect 38344 19184 38350 19236
rect 37458 19156 37464 19168
rect 23400 19128 37464 19156
rect 37458 19116 37464 19128
rect 37516 19116 37522 19168
rect 38010 19156 38016 19168
rect 37971 19128 38016 19156
rect 38010 19116 38016 19128
rect 38068 19116 38074 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1854 18952 1860 18964
rect 1815 18924 1860 18952
rect 1854 18912 1860 18924
rect 1912 18912 1918 18964
rect 2038 18912 2044 18964
rect 2096 18952 2102 18964
rect 2409 18955 2467 18961
rect 2409 18952 2421 18955
rect 2096 18924 2421 18952
rect 2096 18912 2102 18924
rect 2409 18921 2421 18924
rect 2455 18921 2467 18955
rect 2409 18915 2467 18921
rect 20993 18955 21051 18961
rect 20993 18921 21005 18955
rect 21039 18952 21051 18955
rect 21082 18952 21088 18964
rect 21039 18924 21088 18952
rect 21039 18921 21051 18924
rect 20993 18915 21051 18921
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 31754 18912 31760 18964
rect 31812 18952 31818 18964
rect 37277 18955 37335 18961
rect 37277 18952 37289 18955
rect 31812 18924 37289 18952
rect 31812 18912 31818 18924
rect 37277 18921 37289 18924
rect 37323 18921 37335 18955
rect 37277 18915 37335 18921
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 1946 18748 1952 18760
rect 1907 18720 1952 18748
rect 1765 18711 1823 18717
rect 1780 18680 1808 18711
rect 1946 18708 1952 18720
rect 2004 18708 2010 18760
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18748 19763 18751
rect 20070 18748 20076 18760
rect 19751 18720 20076 18748
rect 19751 18717 19763 18720
rect 19705 18711 19763 18717
rect 20070 18708 20076 18720
rect 20128 18708 20134 18760
rect 37292 18748 37320 18915
rect 37829 18751 37887 18757
rect 37829 18748 37841 18751
rect 37292 18720 37841 18748
rect 37829 18717 37841 18720
rect 37875 18717 37887 18751
rect 37829 18711 37887 18717
rect 2314 18680 2320 18692
rect 1780 18652 2320 18680
rect 2314 18640 2320 18652
rect 2372 18640 2378 18692
rect 19889 18683 19947 18689
rect 19889 18649 19901 18683
rect 19935 18680 19947 18683
rect 19935 18652 26234 18680
rect 19935 18649 19947 18652
rect 19889 18643 19947 18649
rect 20346 18612 20352 18624
rect 20307 18584 20352 18612
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 26206 18612 26234 18652
rect 37366 18612 37372 18624
rect 26206 18584 37372 18612
rect 37366 18572 37372 18584
rect 37424 18572 37430 18624
rect 38010 18612 38016 18624
rect 37971 18584 38016 18612
rect 38010 18572 38016 18584
rect 38068 18572 38074 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18272 2102 18284
rect 2685 18275 2743 18281
rect 2685 18272 2697 18275
rect 2096 18244 2697 18272
rect 2096 18232 2102 18244
rect 2685 18241 2697 18244
rect 2731 18241 2743 18275
rect 2685 18235 2743 18241
rect 1596 18176 16574 18204
rect 1596 18145 1624 18176
rect 1581 18139 1639 18145
rect 1581 18105 1593 18139
rect 1627 18105 1639 18139
rect 1581 18099 1639 18105
rect 2225 18139 2283 18145
rect 2225 18105 2237 18139
rect 2271 18136 2283 18139
rect 16546 18136 16574 18176
rect 17954 18136 17960 18148
rect 2271 18108 6914 18136
rect 16546 18108 17960 18136
rect 2271 18105 2283 18108
rect 2225 18099 2283 18105
rect 6886 18068 6914 18108
rect 17954 18096 17960 18108
rect 18012 18096 18018 18148
rect 20714 18136 20720 18148
rect 19168 18108 20720 18136
rect 19168 18068 19196 18108
rect 20714 18096 20720 18108
rect 20772 18096 20778 18148
rect 6886 18040 19196 18068
rect 19521 18071 19579 18077
rect 19521 18037 19533 18071
rect 19567 18068 19579 18071
rect 20070 18068 20076 18080
rect 19567 18040 20076 18068
rect 19567 18037 19579 18040
rect 19521 18031 19579 18037
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1581 17867 1639 17873
rect 1581 17833 1593 17867
rect 1627 17864 1639 17867
rect 1946 17864 1952 17876
rect 1627 17836 1952 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 1394 17756 1400 17808
rect 1452 17796 1458 17808
rect 2041 17799 2099 17805
rect 2041 17796 2053 17799
rect 1452 17768 2053 17796
rect 1452 17756 1458 17768
rect 2041 17765 2053 17768
rect 2087 17765 2099 17799
rect 2041 17759 2099 17765
rect 19889 17731 19947 17737
rect 19889 17697 19901 17731
rect 19935 17728 19947 17731
rect 19935 17700 26234 17728
rect 19935 17697 19947 17700
rect 19889 17691 19947 17697
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17660 1455 17663
rect 1486 17660 1492 17672
rect 1443 17632 1492 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 1486 17620 1492 17632
rect 1544 17620 1550 17672
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 17920 17632 20361 17660
rect 17920 17620 17926 17632
rect 20349 17629 20361 17632
rect 20395 17660 20407 17663
rect 20993 17663 21051 17669
rect 20993 17660 21005 17663
rect 20395 17632 21005 17660
rect 20395 17629 20407 17632
rect 20349 17623 20407 17629
rect 20993 17629 21005 17632
rect 21039 17629 21051 17663
rect 20993 17623 21051 17629
rect 19705 17595 19763 17601
rect 19705 17561 19717 17595
rect 19751 17561 19763 17595
rect 26206 17592 26234 17700
rect 27522 17620 27528 17672
rect 27580 17660 27586 17672
rect 37277 17663 37335 17669
rect 37277 17660 37289 17663
rect 27580 17632 37289 17660
rect 27580 17620 27586 17632
rect 37277 17629 37289 17632
rect 37323 17660 37335 17663
rect 37829 17663 37887 17669
rect 37829 17660 37841 17663
rect 37323 17632 37841 17660
rect 37323 17629 37335 17632
rect 37277 17623 37335 17629
rect 37829 17629 37841 17632
rect 37875 17629 37887 17663
rect 37829 17623 37887 17629
rect 38194 17592 38200 17604
rect 19705 17555 19763 17561
rect 20548 17564 23428 17592
rect 26206 17564 38200 17592
rect 18598 17524 18604 17536
rect 18559 17496 18604 17524
rect 18598 17484 18604 17496
rect 18656 17524 18662 17536
rect 19720 17524 19748 17555
rect 20548 17533 20576 17564
rect 18656 17496 19748 17524
rect 20533 17527 20591 17533
rect 18656 17484 18662 17496
rect 20533 17493 20545 17527
rect 20579 17493 20591 17527
rect 23400 17524 23428 17564
rect 38194 17552 38200 17564
rect 38252 17552 38258 17604
rect 31018 17524 31024 17536
rect 23400 17496 31024 17524
rect 20533 17487 20591 17493
rect 31018 17484 31024 17496
rect 31076 17484 31082 17536
rect 38010 17524 38016 17536
rect 37971 17496 38016 17524
rect 38010 17484 38016 17496
rect 38068 17484 38074 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1486 17280 1492 17332
rect 1544 17320 1550 17332
rect 2041 17323 2099 17329
rect 2041 17320 2053 17323
rect 1544 17292 2053 17320
rect 1544 17280 1550 17292
rect 2041 17289 2053 17292
rect 2087 17289 2099 17323
rect 2041 17283 2099 17289
rect 13906 17212 13912 17264
rect 13964 17252 13970 17264
rect 20349 17255 20407 17261
rect 20349 17252 20361 17255
rect 13964 17224 20361 17252
rect 13964 17212 13970 17224
rect 20349 17221 20361 17224
rect 20395 17252 20407 17255
rect 20993 17255 21051 17261
rect 20993 17252 21005 17255
rect 20395 17224 21005 17252
rect 20395 17221 20407 17224
rect 20349 17215 20407 17221
rect 20993 17221 21005 17224
rect 21039 17221 21051 17255
rect 20993 17215 21051 17221
rect 1394 17184 1400 17196
rect 1355 17156 1400 17184
rect 1394 17144 1400 17156
rect 1452 17184 1458 17196
rect 2593 17187 2651 17193
rect 2593 17184 2605 17187
rect 1452 17156 2605 17184
rect 1452 17144 1458 17156
rect 2593 17153 2605 17156
rect 2639 17153 2651 17187
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 2593 17147 2651 17153
rect 18984 17156 19625 17184
rect 1581 17051 1639 17057
rect 1581 17017 1593 17051
rect 1627 17048 1639 17051
rect 18598 17048 18604 17060
rect 1627 17020 18604 17048
rect 1627 17017 1639 17020
rect 1581 17011 1639 17017
rect 18598 17008 18604 17020
rect 18656 17008 18662 17060
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 18984 16989 19012 17156
rect 19613 17153 19625 17156
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 31018 17144 31024 17196
rect 31076 17184 31082 17196
rect 37829 17187 37887 17193
rect 37829 17184 37841 17187
rect 31076 17156 37841 17184
rect 31076 17144 31082 17156
rect 37829 17153 37841 17156
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17116 20591 17119
rect 20579 17088 35894 17116
rect 20579 17085 20591 17088
rect 20533 17079 20591 17085
rect 19797 17051 19855 17057
rect 19797 17017 19809 17051
rect 19843 17048 19855 17051
rect 35866 17048 35894 17088
rect 38102 17048 38108 17060
rect 19843 17020 26234 17048
rect 35866 17020 38108 17048
rect 19843 17017 19855 17020
rect 19797 17011 19855 17017
rect 18969 16983 19027 16989
rect 18969 16980 18981 16983
rect 15160 16952 18981 16980
rect 15160 16940 15166 16952
rect 18969 16949 18981 16952
rect 19015 16949 19027 16983
rect 26206 16980 26234 17020
rect 38102 17008 38108 17020
rect 38160 17008 38166 17060
rect 37734 16980 37740 16992
rect 26206 16952 37740 16980
rect 18969 16943 19027 16949
rect 37734 16940 37740 16952
rect 37792 16940 37798 16992
rect 38010 16980 38016 16992
rect 37971 16952 38016 16980
rect 38010 16940 38016 16952
rect 38068 16940 38074 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 20714 16776 20720 16788
rect 20675 16748 20720 16776
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 20732 16640 20760 16736
rect 20088 16612 20760 16640
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16572 1455 16575
rect 1486 16572 1492 16584
rect 1443 16544 1492 16572
rect 1443 16541 1455 16544
rect 1397 16535 1455 16541
rect 1486 16532 1492 16544
rect 1544 16532 1550 16584
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16572 2102 16584
rect 2685 16575 2743 16581
rect 2685 16572 2697 16575
rect 2096 16544 2697 16572
rect 2096 16532 2102 16544
rect 2685 16541 2697 16544
rect 2731 16541 2743 16575
rect 2685 16535 2743 16541
rect 17954 16532 17960 16584
rect 18012 16572 18018 16584
rect 19242 16572 19248 16584
rect 18012 16544 19248 16572
rect 18012 16532 18018 16544
rect 19242 16532 19248 16544
rect 19300 16572 19306 16584
rect 20088 16581 20116 16612
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 19300 16544 19441 16572
rect 19300 16532 19306 16544
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16574 20131 16575
rect 37829 16575 37887 16581
rect 20119 16546 20153 16574
rect 20119 16541 20131 16546
rect 20073 16535 20131 16541
rect 37829 16541 37841 16575
rect 37875 16541 37887 16575
rect 37829 16535 37887 16541
rect 37277 16507 37335 16513
rect 37277 16504 37289 16507
rect 19628 16476 37289 16504
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 2222 16436 2228 16448
rect 2183 16408 2228 16436
rect 2222 16396 2228 16408
rect 2280 16396 2286 16448
rect 19628 16445 19656 16476
rect 37277 16473 37289 16476
rect 37323 16504 37335 16507
rect 37844 16504 37872 16535
rect 37323 16476 37872 16504
rect 37323 16473 37335 16476
rect 37277 16467 37335 16473
rect 19613 16439 19671 16445
rect 19613 16405 19625 16439
rect 19659 16405 19671 16439
rect 19613 16399 19671 16405
rect 20257 16439 20315 16445
rect 20257 16405 20269 16439
rect 20303 16436 20315 16439
rect 37182 16436 37188 16448
rect 20303 16408 37188 16436
rect 20303 16405 20315 16408
rect 20257 16399 20315 16405
rect 37182 16396 37188 16408
rect 37240 16396 37246 16448
rect 38010 16436 38016 16448
rect 37971 16408 38016 16436
rect 38010 16396 38016 16408
rect 38068 16396 38074 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 1636 16204 6914 16232
rect 1636 16192 1642 16204
rect 1486 16124 1492 16176
rect 1544 16164 1550 16176
rect 2041 16167 2099 16173
rect 2041 16164 2053 16167
rect 1544 16136 2053 16164
rect 1544 16124 1550 16136
rect 2041 16133 2053 16136
rect 2087 16133 2099 16167
rect 2041 16127 2099 16133
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 6886 16096 6914 16204
rect 19242 16192 19248 16244
rect 19300 16232 19306 16244
rect 19337 16235 19395 16241
rect 19337 16232 19349 16235
rect 19300 16204 19349 16232
rect 19300 16192 19306 16204
rect 19337 16201 19349 16204
rect 19383 16201 19395 16235
rect 19337 16195 19395 16201
rect 37182 16192 37188 16244
rect 37240 16232 37246 16244
rect 37277 16235 37335 16241
rect 37277 16232 37289 16235
rect 37240 16204 37289 16232
rect 37240 16192 37246 16204
rect 37277 16201 37289 16204
rect 37323 16201 37335 16235
rect 37277 16195 37335 16201
rect 19797 16099 19855 16105
rect 19797 16096 19809 16099
rect 6886 16068 19809 16096
rect 19797 16065 19809 16068
rect 19843 16096 19855 16099
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 19843 16068 20453 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 37292 16096 37320 16195
rect 37829 16099 37887 16105
rect 37829 16096 37841 16099
rect 37292 16068 37841 16096
rect 20441 16059 20499 16065
rect 37829 16065 37841 16068
rect 37875 16065 37887 16099
rect 37829 16059 37887 16065
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 15102 15960 15108 15972
rect 1627 15932 15108 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 15102 15920 15108 15932
rect 15160 15920 15166 15972
rect 19981 15963 20039 15969
rect 19981 15929 19993 15963
rect 20027 15960 20039 15963
rect 33134 15960 33140 15972
rect 20027 15932 33140 15960
rect 20027 15929 20039 15932
rect 19981 15923 20039 15929
rect 33134 15920 33140 15932
rect 33192 15920 33198 15972
rect 38010 15892 38016 15904
rect 37971 15864 38016 15892
rect 38010 15852 38016 15864
rect 38068 15852 38074 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1486 15648 1492 15700
rect 1544 15688 1550 15700
rect 2041 15691 2099 15697
rect 2041 15688 2053 15691
rect 1544 15660 2053 15688
rect 1544 15648 1550 15660
rect 2041 15657 2053 15660
rect 2087 15657 2099 15691
rect 2041 15651 2099 15657
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15484 1458 15496
rect 2593 15487 2651 15493
rect 2593 15484 2605 15487
rect 1452 15456 2605 15484
rect 1452 15444 1458 15456
rect 2593 15453 2605 15456
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 13906 15416 13912 15428
rect 1596 15388 13912 15416
rect 1596 15357 1624 15388
rect 13906 15376 13912 15388
rect 13964 15376 13970 15428
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 33134 15104 33140 15156
rect 33192 15144 33198 15156
rect 37277 15147 37335 15153
rect 37277 15144 37289 15147
rect 33192 15116 37289 15144
rect 33192 15104 33198 15116
rect 37277 15113 37289 15116
rect 37323 15113 37335 15147
rect 37277 15107 37335 15113
rect 2222 15036 2228 15088
rect 2280 15076 2286 15088
rect 2280 15048 6914 15076
rect 2280 15036 2286 15048
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 2038 15008 2044 15020
rect 1999 14980 2044 15008
rect 2038 14968 2044 14980
rect 2096 15008 2102 15020
rect 2685 15011 2743 15017
rect 2685 15008 2697 15011
rect 2096 14980 2697 15008
rect 2096 14968 2102 14980
rect 2685 14977 2697 14980
rect 2731 14977 2743 15011
rect 6886 15008 6914 15048
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 6886 14980 19993 15008
rect 2685 14971 2743 14977
rect 19981 14977 19993 14980
rect 20027 15008 20039 15011
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 20027 14980 20637 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 37292 15008 37320 15107
rect 37829 15011 37887 15017
rect 37829 15008 37841 15011
rect 37292 14980 37841 15008
rect 20625 14971 20683 14977
rect 37829 14977 37841 14980
rect 37875 14977 37887 15011
rect 37829 14971 37887 14977
rect 37274 14940 37280 14952
rect 1596 14912 16574 14940
rect 1596 14881 1624 14912
rect 1581 14875 1639 14881
rect 1581 14841 1593 14875
rect 1627 14841 1639 14875
rect 1581 14835 1639 14841
rect 2225 14875 2283 14881
rect 2225 14841 2237 14875
rect 2271 14872 2283 14875
rect 16546 14872 16574 14912
rect 26206 14912 37280 14940
rect 19978 14872 19984 14884
rect 2271 14844 6914 14872
rect 16546 14844 19984 14872
rect 2271 14841 2283 14844
rect 2225 14835 2283 14841
rect 6886 14804 6914 14844
rect 19978 14832 19984 14844
rect 20036 14832 20042 14884
rect 20165 14875 20223 14881
rect 20165 14841 20177 14875
rect 20211 14872 20223 14875
rect 26206 14872 26234 14912
rect 37274 14900 37280 14912
rect 37332 14900 37338 14952
rect 38010 14872 38016 14884
rect 20211 14844 26234 14872
rect 37971 14844 38016 14872
rect 20211 14841 20223 14844
rect 20165 14835 20223 14841
rect 38010 14832 38016 14844
rect 38068 14832 38074 14884
rect 19426 14804 19432 14816
rect 6886 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1486 14560 1492 14612
rect 1544 14600 1550 14612
rect 2041 14603 2099 14609
rect 2041 14600 2053 14603
rect 1544 14572 2053 14600
rect 1544 14560 1550 14572
rect 2041 14569 2053 14572
rect 2087 14569 2099 14603
rect 37274 14600 37280 14612
rect 37235 14572 37280 14600
rect 2041 14563 2099 14569
rect 37274 14560 37280 14572
rect 37332 14560 37338 14612
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14396 1458 14408
rect 2593 14399 2651 14405
rect 2593 14396 2605 14399
rect 1452 14368 2605 14396
rect 1452 14356 1458 14368
rect 2593 14365 2605 14368
rect 2639 14365 2651 14399
rect 19978 14396 19984 14408
rect 19939 14368 19984 14396
rect 2593 14359 2651 14365
rect 19978 14356 19984 14368
rect 20036 14396 20042 14408
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 20036 14368 20637 14396
rect 20036 14356 20042 14368
rect 20625 14365 20637 14368
rect 20671 14365 20683 14399
rect 37292 14396 37320 14560
rect 37829 14399 37887 14405
rect 37829 14396 37841 14399
rect 37292 14368 37841 14396
rect 20625 14359 20683 14365
rect 37829 14365 37841 14368
rect 37875 14365 37887 14399
rect 37829 14359 37887 14365
rect 20180 14300 26234 14328
rect 1578 14260 1584 14272
rect 1539 14232 1584 14260
rect 1578 14220 1584 14232
rect 1636 14220 1642 14272
rect 20180 14269 20208 14300
rect 20165 14263 20223 14269
rect 20165 14229 20177 14263
rect 20211 14229 20223 14263
rect 26206 14260 26234 14300
rect 37182 14260 37188 14272
rect 26206 14232 37188 14260
rect 20165 14223 20223 14229
rect 37182 14220 37188 14232
rect 37240 14220 37246 14272
rect 38010 14260 38016 14272
rect 37971 14232 38016 14260
rect 38010 14220 38016 14232
rect 38068 14220 38074 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1627 14028 6914 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 6886 13988 6914 14028
rect 37182 14016 37188 14068
rect 37240 14056 37246 14068
rect 37277 14059 37335 14065
rect 37277 14056 37289 14059
rect 37240 14028 37289 14056
rect 37240 14016 37246 14028
rect 37277 14025 37289 14028
rect 37323 14025 37335 14059
rect 37277 14019 37335 14025
rect 20346 13988 20352 14000
rect 6886 13960 20352 13988
rect 20346 13948 20352 13960
rect 20404 13948 20410 14000
rect 1394 13920 1400 13932
rect 1355 13892 1400 13920
rect 1394 13880 1400 13892
rect 1452 13880 1458 13932
rect 2038 13920 2044 13932
rect 1999 13892 2044 13920
rect 2038 13880 2044 13892
rect 2096 13920 2102 13932
rect 2685 13923 2743 13929
rect 2685 13920 2697 13923
rect 2096 13892 2697 13920
rect 2096 13880 2102 13892
rect 2685 13889 2697 13892
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 19484 13892 19993 13920
rect 19484 13880 19490 13892
rect 19981 13889 19993 13892
rect 20027 13920 20039 13923
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20027 13892 20637 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 37292 13920 37320 14019
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 37292 13892 37841 13920
rect 20625 13883 20683 13889
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 1412 13852 1440 13880
rect 3237 13855 3295 13861
rect 3237 13852 3249 13855
rect 1412 13824 3249 13852
rect 3237 13821 3249 13824
rect 3283 13821 3295 13855
rect 37182 13852 37188 13864
rect 3237 13815 3295 13821
rect 20180 13824 37188 13852
rect 20180 13793 20208 13824
rect 37182 13812 37188 13824
rect 37240 13812 37246 13864
rect 20165 13787 20223 13793
rect 20165 13753 20177 13787
rect 20211 13753 20223 13787
rect 20165 13747 20223 13753
rect 2222 13716 2228 13728
rect 2183 13688 2228 13716
rect 2222 13676 2228 13688
rect 2280 13676 2286 13728
rect 38010 13716 38016 13728
rect 37971 13688 38016 13716
rect 38010 13676 38016 13688
rect 38068 13676 38074 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 37182 13472 37188 13524
rect 37240 13512 37246 13524
rect 37277 13515 37335 13521
rect 37277 13512 37289 13515
rect 37240 13484 37289 13512
rect 37240 13472 37246 13484
rect 37277 13481 37289 13484
rect 37323 13481 37335 13515
rect 37277 13475 37335 13481
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 19334 13376 19340 13388
rect 1995 13348 19340 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 2225 13311 2283 13317
rect 2225 13308 2237 13311
rect 2188 13280 2237 13308
rect 2188 13268 2194 13280
rect 2225 13277 2237 13280
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13308 2743 13311
rect 2774 13308 2780 13320
rect 2731 13280 2780 13308
rect 2731 13277 2743 13280
rect 2685 13271 2743 13277
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 37292 13308 37320 13475
rect 37829 13311 37887 13317
rect 37829 13308 37841 13311
rect 37292 13280 37841 13308
rect 37829 13277 37841 13280
rect 37875 13277 37887 13311
rect 37829 13271 37887 13277
rect 2869 13175 2927 13181
rect 2869 13141 2881 13175
rect 2915 13172 2927 13175
rect 15194 13172 15200 13184
rect 2915 13144 15200 13172
rect 2915 13141 2927 13144
rect 2869 13135 2927 13141
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 38010 13172 38016 13184
rect 37971 13144 38016 13172
rect 38010 13132 38016 13144
rect 38068 13132 38074 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 2222 12928 2228 12980
rect 2280 12968 2286 12980
rect 2280 12940 16574 12968
rect 2280 12928 2286 12940
rect 2774 12900 2780 12912
rect 2735 12872 2780 12900
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 16546 12832 16574 12940
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 1995 12804 6914 12832
rect 16546 12804 19809 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2222 12764 2228 12776
rect 2183 12736 2228 12764
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 6886 12764 6914 12804
rect 19797 12801 19809 12804
rect 19843 12832 19855 12835
rect 20441 12835 20499 12841
rect 20441 12832 20453 12835
rect 19843 12804 20453 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 20441 12801 20453 12804
rect 20487 12801 20499 12835
rect 20441 12795 20499 12801
rect 18414 12764 18420 12776
rect 6886 12736 18420 12764
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 19981 12699 20039 12705
rect 19981 12665 19993 12699
rect 20027 12696 20039 12699
rect 20027 12668 26234 12696
rect 20027 12665 20039 12668
rect 19981 12659 20039 12665
rect 26206 12628 26234 12668
rect 36998 12628 37004 12640
rect 26206 12600 37004 12628
rect 36998 12588 37004 12600
rect 37056 12588 37062 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 2130 12424 2136 12436
rect 2091 12396 2136 12424
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 2222 12384 2228 12436
rect 2280 12424 2286 12436
rect 2593 12427 2651 12433
rect 2593 12424 2605 12427
rect 2280 12396 2605 12424
rect 2280 12384 2286 12396
rect 2593 12393 2605 12396
rect 2639 12393 2651 12427
rect 2593 12387 2651 12393
rect 36998 12384 37004 12436
rect 37056 12424 37062 12436
rect 37277 12427 37335 12433
rect 37277 12424 37289 12427
rect 37056 12396 37289 12424
rect 37056 12384 37062 12396
rect 37277 12393 37289 12396
rect 37323 12393 37335 12427
rect 37277 12387 37335 12393
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 15252 12192 19809 12220
rect 15252 12180 15258 12192
rect 19797 12189 19809 12192
rect 19843 12220 19855 12223
rect 20441 12223 20499 12229
rect 20441 12220 20453 12223
rect 19843 12192 20453 12220
rect 19843 12189 19855 12192
rect 19797 12183 19855 12189
rect 20441 12189 20453 12192
rect 20487 12189 20499 12223
rect 37292 12220 37320 12387
rect 37829 12223 37887 12229
rect 37829 12220 37841 12223
rect 37292 12192 37841 12220
rect 20441 12183 20499 12189
rect 37829 12189 37841 12192
rect 37875 12189 37887 12223
rect 37829 12183 37887 12189
rect 15286 12152 15292 12164
rect 1596 12124 15292 12152
rect 1596 12093 1624 12124
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 19996 12124 26234 12152
rect 19996 12093 20024 12124
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12053 1639 12087
rect 1581 12047 1639 12053
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12053 20039 12087
rect 26206 12084 26234 12124
rect 37182 12084 37188 12096
rect 26206 12056 37188 12084
rect 19981 12047 20039 12053
rect 37182 12044 37188 12056
rect 37240 12044 37246 12096
rect 38010 12084 38016 12096
rect 37971 12056 38016 12084
rect 38010 12044 38016 12056
rect 38068 12044 38074 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 37182 11840 37188 11892
rect 37240 11880 37246 11892
rect 37277 11883 37335 11889
rect 37277 11880 37289 11883
rect 37240 11852 37289 11880
rect 37240 11840 37246 11852
rect 37277 11849 37289 11852
rect 37323 11849 37335 11883
rect 37277 11843 37335 11849
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 14458 11744 14464 11756
rect 1995 11716 14464 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 37292 11744 37320 11843
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 37292 11716 37841 11744
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11676 2286 11688
rect 2685 11679 2743 11685
rect 2685 11676 2697 11679
rect 2280 11648 2697 11676
rect 2280 11636 2286 11648
rect 2685 11645 2697 11648
rect 2731 11645 2743 11679
rect 2685 11639 2743 11645
rect 38010 11540 38016 11552
rect 37971 11512 38016 11540
rect 38010 11500 38016 11512
rect 38068 11500 38074 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1486 11296 1492 11348
rect 1544 11336 1550 11348
rect 2041 11339 2099 11345
rect 2041 11336 2053 11339
rect 1544 11308 2053 11336
rect 1544 11296 1550 11308
rect 2041 11305 2053 11308
rect 2087 11305 2099 11339
rect 2041 11299 2099 11305
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 19981 11271 20039 11277
rect 1627 11240 6914 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11132 1458 11144
rect 2593 11135 2651 11141
rect 2593 11132 2605 11135
rect 1452 11104 2605 11132
rect 1452 11092 1458 11104
rect 2593 11101 2605 11104
rect 2639 11101 2651 11135
rect 6886 11132 6914 11240
rect 19981 11237 19993 11271
rect 20027 11268 20039 11271
rect 38010 11268 38016 11280
rect 20027 11240 26234 11268
rect 37971 11240 38016 11268
rect 20027 11237 20039 11240
rect 19981 11231 20039 11237
rect 19797 11135 19855 11141
rect 19797 11132 19809 11135
rect 6886 11104 19809 11132
rect 2593 11095 2651 11101
rect 19797 11101 19809 11104
rect 19843 11132 19855 11135
rect 20441 11135 20499 11141
rect 20441 11132 20453 11135
rect 19843 11104 20453 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 20441 11101 20453 11104
rect 20487 11101 20499 11135
rect 26206 11132 26234 11240
rect 38010 11228 38016 11240
rect 38068 11228 38074 11280
rect 37829 11135 37887 11141
rect 37829 11132 37841 11135
rect 26206 11104 37841 11132
rect 20441 11095 20499 11101
rect 37829 11101 37841 11104
rect 37875 11101 37887 11135
rect 37829 11095 37887 11101
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10656 2102 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2096 10628 2697 10656
rect 2096 10616 2102 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 37829 10659 37887 10665
rect 37829 10656 37841 10659
rect 2685 10619 2743 10625
rect 37292 10628 37841 10656
rect 2225 10523 2283 10529
rect 2225 10489 2237 10523
rect 2271 10520 2283 10523
rect 19702 10520 19708 10532
rect 2271 10492 19708 10520
rect 2271 10489 2283 10492
rect 2225 10483 2283 10489
rect 19702 10480 19708 10492
rect 19760 10480 19766 10532
rect 37292 10464 37320 10628
rect 37829 10625 37841 10628
rect 37875 10625 37887 10659
rect 37829 10619 37887 10625
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 37274 10452 37280 10464
rect 37235 10424 37280 10452
rect 37274 10412 37280 10424
rect 37332 10412 37338 10464
rect 38010 10452 38016 10464
rect 37971 10424 38016 10452
rect 38010 10412 38016 10424
rect 38068 10412 38074 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 13814 10248 13820 10260
rect 1636 10220 13820 10248
rect 1636 10208 1642 10220
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 1995 10084 6914 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 2222 10044 2228 10056
rect 2183 10016 2228 10044
rect 2222 10004 2228 10016
rect 2280 10044 2286 10056
rect 2685 10047 2743 10053
rect 2685 10044 2697 10047
rect 2280 10016 2697 10044
rect 2280 10004 2286 10016
rect 2685 10013 2697 10016
rect 2731 10013 2743 10047
rect 6886 10044 6914 10084
rect 18506 10044 18512 10056
rect 6886 10016 18512 10044
rect 2685 10007 2743 10013
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 19702 10044 19708 10056
rect 19663 10016 19708 10044
rect 19702 10004 19708 10016
rect 19760 10044 19766 10056
rect 20349 10047 20407 10053
rect 20349 10044 20361 10047
rect 19760 10016 20361 10044
rect 19760 10004 19766 10016
rect 20349 10013 20361 10016
rect 20395 10013 20407 10047
rect 20349 10007 20407 10013
rect 19904 9948 26234 9976
rect 19904 9917 19932 9948
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9877 19947 9911
rect 26206 9908 26234 9948
rect 37274 9908 37280 9920
rect 26206 9880 37280 9908
rect 19889 9871 19947 9877
rect 37274 9868 37280 9880
rect 37332 9868 37338 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2041 9707 2099 9713
rect 2041 9704 2053 9707
rect 1452 9676 2053 9704
rect 1452 9664 1458 9676
rect 2041 9673 2053 9676
rect 2087 9673 2099 9707
rect 2041 9667 2099 9673
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 19702 9568 19708 9580
rect 19663 9540 19708 9568
rect 19702 9528 19708 9540
rect 19760 9568 19766 9580
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 19760 9540 20361 9568
rect 19760 9528 19766 9540
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 37829 9571 37887 9577
rect 37829 9568 37841 9571
rect 20349 9531 20407 9537
rect 26206 9540 37841 9568
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 19889 9435 19947 9441
rect 1627 9404 6914 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 6886 9364 6914 9404
rect 19889 9401 19901 9435
rect 19935 9432 19947 9435
rect 26206 9432 26234 9540
rect 37829 9537 37841 9540
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 38010 9432 38016 9444
rect 19935 9404 26234 9432
rect 37971 9404 38016 9432
rect 19935 9401 19947 9404
rect 19889 9395 19947 9401
rect 38010 9392 38016 9404
rect 38068 9392 38074 9444
rect 18414 9364 18420 9376
rect 6886 9336 18420 9364
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 2041 9163 2099 9169
rect 2041 9160 2053 9163
rect 1544 9132 2053 9160
rect 1544 9120 1550 9132
rect 2041 9129 2053 9132
rect 2087 9129 2099 9163
rect 2041 9123 2099 9129
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 1627 9064 6914 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8956 1458 8968
rect 2593 8959 2651 8965
rect 2593 8956 2605 8959
rect 1452 8928 2605 8956
rect 1452 8916 1458 8928
rect 2593 8925 2605 8928
rect 2639 8925 2651 8959
rect 6886 8956 6914 9064
rect 19702 8956 19708 8968
rect 6886 8928 19708 8956
rect 2593 8919 2651 8925
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 37829 8959 37887 8965
rect 37829 8956 37841 8959
rect 37292 8928 37841 8956
rect 13814 8848 13820 8900
rect 13872 8888 13878 8900
rect 20257 8891 20315 8897
rect 20257 8888 20269 8891
rect 13872 8860 20269 8888
rect 13872 8848 13878 8860
rect 20257 8857 20269 8860
rect 20303 8888 20315 8891
rect 20622 8888 20628 8900
rect 20303 8860 20628 8888
rect 20303 8857 20315 8860
rect 20257 8851 20315 8857
rect 20622 8848 20628 8860
rect 20680 8848 20686 8900
rect 37292 8832 37320 8928
rect 37829 8925 37841 8928
rect 37875 8925 37887 8959
rect 37829 8919 37887 8925
rect 19337 8823 19395 8829
rect 19337 8789 19349 8823
rect 19383 8820 19395 8823
rect 19426 8820 19432 8832
rect 19383 8792 19432 8820
rect 19383 8789 19395 8792
rect 19337 8783 19395 8789
rect 19426 8780 19432 8792
rect 19484 8820 19490 8832
rect 20809 8823 20867 8829
rect 20809 8820 20821 8823
rect 19484 8792 20821 8820
rect 19484 8780 19490 8792
rect 20809 8789 20821 8792
rect 20855 8789 20867 8823
rect 37274 8820 37280 8832
rect 37235 8792 37280 8820
rect 20809 8783 20867 8789
rect 37274 8780 37280 8792
rect 37332 8780 37338 8832
rect 38010 8820 38016 8832
rect 37971 8792 38016 8820
rect 38010 8780 38016 8792
rect 38068 8780 38074 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 15286 8576 15292 8628
rect 15344 8616 15350 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 15344 8588 19073 8616
rect 15344 8576 15350 8588
rect 19061 8585 19073 8588
rect 19107 8616 19119 8619
rect 19107 8588 19196 8616
rect 19107 8585 19119 8588
rect 19061 8579 19119 8585
rect 2314 8548 2320 8560
rect 2275 8520 2320 8548
rect 2314 8508 2320 8520
rect 2372 8508 2378 8560
rect 2501 8551 2559 8557
rect 2501 8517 2513 8551
rect 2547 8548 2559 8551
rect 2547 8520 19012 8548
rect 2547 8517 2559 8520
rect 2501 8511 2559 8517
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 18598 8412 18604 8424
rect 6886 8384 18604 8412
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 6886 8344 6914 8384
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 1627 8316 6914 8344
rect 18984 8344 19012 8520
rect 19168 8480 19196 8588
rect 37274 8548 37280 8560
rect 26206 8520 37280 8548
rect 19797 8483 19855 8489
rect 19797 8480 19809 8483
rect 19168 8452 19809 8480
rect 19797 8449 19809 8452
rect 19843 8449 19855 8483
rect 20622 8480 20628 8492
rect 20583 8452 20628 8480
rect 19797 8443 19855 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 19613 8415 19671 8421
rect 19613 8412 19625 8415
rect 19484 8384 19625 8412
rect 19484 8372 19490 8384
rect 19613 8381 19625 8384
rect 19659 8412 19671 8415
rect 20441 8415 20499 8421
rect 20441 8412 20453 8415
rect 19659 8384 20453 8412
rect 19659 8381 19671 8384
rect 19613 8375 19671 8381
rect 20441 8381 20453 8384
rect 20487 8381 20499 8415
rect 20441 8375 20499 8381
rect 26206 8344 26234 8520
rect 37274 8508 37280 8520
rect 37332 8508 37338 8560
rect 37366 8440 37372 8492
rect 37424 8480 37430 8492
rect 37829 8483 37887 8489
rect 37829 8480 37841 8483
rect 37424 8452 37841 8480
rect 37424 8440 37430 8452
rect 37829 8449 37841 8452
rect 37875 8449 37887 8483
rect 37829 8443 37887 8449
rect 38010 8344 38016 8356
rect 18984 8316 26234 8344
rect 37971 8316 38016 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 38010 8304 38016 8316
rect 38068 8304 38074 8356
rect 19981 8279 20039 8285
rect 19981 8245 19993 8279
rect 20027 8276 20039 8279
rect 20622 8276 20628 8288
rect 20027 8248 20628 8276
rect 20027 8245 20039 8248
rect 19981 8239 20039 8245
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 20809 8279 20867 8285
rect 20809 8245 20821 8279
rect 20855 8276 20867 8279
rect 21266 8276 21272 8288
rect 20855 8248 21272 8276
rect 20855 8245 20867 8248
rect 20809 8239 20867 8245
rect 21266 8236 21272 8248
rect 21324 8236 21330 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 2041 8075 2099 8081
rect 2041 8072 2053 8075
rect 1452 8044 2053 8072
rect 1452 8032 1458 8044
rect 2041 8041 2053 8044
rect 2087 8041 2099 8075
rect 2041 8035 2099 8041
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 18472 8044 18613 8072
rect 18472 8032 18478 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 2314 8004 2320 8016
rect 1627 7976 2320 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 18616 7936 18644 8035
rect 18616 7908 19840 7936
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7868 1458 7880
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 1452 7840 2605 7868
rect 1452 7828 1458 7840
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 19426 7828 19432 7880
rect 19484 7868 19490 7880
rect 19812 7877 19840 7908
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19484 7840 19625 7868
rect 19484 7828 19490 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7837 19855 7871
rect 20622 7868 20628 7880
rect 20583 7840 20628 7868
rect 19797 7831 19855 7837
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 21266 7868 21272 7880
rect 21227 7840 21272 7868
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 37829 7871 37887 7877
rect 37829 7837 37841 7871
rect 37875 7837 37887 7871
rect 37829 7831 37887 7837
rect 37366 7800 37372 7812
rect 20824 7772 37372 7800
rect 19981 7735 20039 7741
rect 19981 7701 19993 7735
rect 20027 7732 20039 7735
rect 20622 7732 20628 7744
rect 20027 7704 20628 7732
rect 20027 7701 20039 7704
rect 19981 7695 20039 7701
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 20824 7741 20852 7772
rect 37366 7760 37372 7772
rect 37424 7760 37430 7812
rect 20809 7735 20867 7741
rect 20809 7701 20821 7735
rect 20855 7701 20867 7735
rect 20809 7695 20867 7701
rect 21453 7735 21511 7741
rect 21453 7701 21465 7735
rect 21499 7732 21511 7735
rect 37844 7732 37872 7831
rect 38010 7732 38016 7744
rect 21499 7704 37872 7732
rect 37971 7704 38016 7732
rect 21499 7701 21511 7704
rect 21453 7695 21511 7701
rect 38010 7692 38016 7704
rect 38068 7692 38074 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 18598 7528 18604 7540
rect 18559 7500 18604 7528
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 1762 7352 1768 7404
rect 1820 7392 1826 7404
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1820 7364 1869 7392
rect 1820 7352 1826 7364
rect 1857 7361 1869 7364
rect 1903 7392 1915 7395
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 1903 7364 2513 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 18616 7392 18644 7488
rect 19153 7395 19211 7401
rect 19153 7392 19165 7395
rect 18616 7364 19165 7392
rect 2501 7355 2559 7361
rect 19153 7361 19165 7364
rect 19199 7361 19211 7395
rect 19153 7355 19211 7361
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 19426 7392 19432 7404
rect 19383 7364 19432 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 19352 7324 19380 7355
rect 19426 7352 19432 7364
rect 19484 7392 19490 7404
rect 19981 7395 20039 7401
rect 19981 7392 19993 7395
rect 19484 7364 19993 7392
rect 19484 7352 19490 7364
rect 19981 7361 19993 7364
rect 20027 7392 20039 7395
rect 20070 7392 20076 7404
rect 20027 7364 20076 7392
rect 20027 7361 20039 7364
rect 19981 7355 20039 7361
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20622 7392 20628 7404
rect 20583 7364 20628 7392
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 18064 7296 19380 7324
rect 18064 7265 18092 7296
rect 2041 7259 2099 7265
rect 2041 7225 2053 7259
rect 2087 7256 2099 7259
rect 18049 7259 18107 7265
rect 18049 7256 18061 7259
rect 2087 7228 18061 7256
rect 2087 7225 2099 7228
rect 2041 7219 2099 7225
rect 18049 7225 18061 7228
rect 18095 7225 18107 7259
rect 18049 7219 18107 7225
rect 19518 7188 19524 7200
rect 19479 7160 19524 7188
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 20809 7191 20867 7197
rect 20809 7157 20821 7191
rect 20855 7188 20867 7191
rect 37826 7188 37832 7200
rect 20855 7160 37832 7188
rect 20855 7157 20867 7160
rect 20809 7151 20867 7157
rect 37826 7148 37832 7160
rect 37884 7148 37890 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1762 6780 1768 6792
rect 1723 6752 1768 6780
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2774 6780 2780 6792
rect 2639 6752 2780 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 1964 6644 1992 6743
rect 2774 6740 2780 6752
rect 2832 6780 2838 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2832 6752 3065 6780
rect 2832 6740 2838 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 20165 6783 20223 6789
rect 20165 6780 20177 6783
rect 19576 6752 20177 6780
rect 19576 6740 19582 6752
rect 20165 6749 20177 6752
rect 20211 6749 20223 6783
rect 37826 6780 37832 6792
rect 37787 6752 37832 6780
rect 20165 6743 20223 6749
rect 37826 6740 37832 6752
rect 37884 6740 37890 6792
rect 2409 6647 2467 6653
rect 2409 6644 2421 6647
rect 1964 6616 2421 6644
rect 2409 6613 2421 6616
rect 2455 6613 2467 6647
rect 2409 6607 2467 6613
rect 20349 6647 20407 6653
rect 20349 6613 20361 6647
rect 20395 6644 20407 6647
rect 37826 6644 37832 6656
rect 20395 6616 37832 6644
rect 20395 6613 20407 6616
rect 20349 6607 20407 6613
rect 37826 6604 37832 6616
rect 37884 6604 37890 6656
rect 38010 6644 38016 6656
rect 37971 6616 38016 6644
rect 38010 6604 38016 6616
rect 38068 6604 38074 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 2130 6304 2136 6316
rect 1719 6276 2136 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 20070 6264 20076 6316
rect 20128 6304 20134 6316
rect 20349 6307 20407 6313
rect 20349 6304 20361 6307
rect 20128 6276 20361 6304
rect 20128 6264 20134 6276
rect 20349 6273 20361 6276
rect 20395 6304 20407 6307
rect 20993 6307 21051 6313
rect 20993 6304 21005 6307
rect 20395 6276 21005 6304
rect 20395 6273 20407 6276
rect 20349 6267 20407 6273
rect 20993 6273 21005 6276
rect 21039 6273 21051 6307
rect 37826 6304 37832 6316
rect 37787 6276 37832 6304
rect 20993 6267 21051 6273
rect 37826 6264 37832 6276
rect 37884 6264 37890 6316
rect 20441 6171 20499 6177
rect 20441 6137 20453 6171
rect 20487 6168 20499 6171
rect 20487 6140 26234 6168
rect 20487 6137 20499 6140
rect 20441 6131 20499 6137
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 26206 6100 26234 6140
rect 37826 6100 37832 6112
rect 26206 6072 37832 6100
rect 37826 6060 37832 6072
rect 37884 6060 37890 6112
rect 38010 6100 38016 6112
rect 37971 6072 38016 6100
rect 38010 6060 38016 6072
rect 38068 6060 38074 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 37826 5692 37832 5704
rect 37787 5664 37832 5692
rect 37826 5652 37832 5664
rect 37884 5652 37890 5704
rect 1394 5584 1400 5636
rect 1452 5624 1458 5636
rect 1489 5627 1547 5633
rect 1489 5624 1501 5627
rect 1452 5596 1501 5624
rect 1452 5584 1458 5596
rect 1489 5593 1501 5596
rect 1535 5593 1547 5627
rect 1489 5587 1547 5593
rect 1946 5584 1952 5636
rect 2004 5624 2010 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 2004 5596 3249 5624
rect 2004 5584 2010 5596
rect 3237 5593 3249 5596
rect 3283 5593 3295 5627
rect 3237 5587 3295 5593
rect 38010 5556 38016 5568
rect 37971 5528 38016 5556
rect 38010 5516 38016 5528
rect 38068 5516 38074 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1762 5352 1768 5364
rect 1627 5324 1768 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 2130 5352 2136 5364
rect 2091 5324 2136 5352
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 2685 5287 2743 5293
rect 2685 5284 2697 5287
rect 1412 5256 2697 5284
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1412 5225 1440 5256
rect 2685 5253 2697 5256
rect 2731 5253 2743 5287
rect 2685 5247 2743 5253
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1360 5188 1409 5216
rect 1360 5176 1366 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1854 5176 1860 5228
rect 1912 5216 1918 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1912 5188 2053 5216
rect 1912 5176 1918 5188
rect 2041 5185 2053 5188
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2774 5216 2780 5228
rect 2271 5188 2780 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 37829 5219 37887 5225
rect 37829 5216 37841 5219
rect 37292 5188 37841 5216
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 37292 5021 37320 5188
rect 37829 5185 37841 5188
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 37277 5015 37335 5021
rect 37277 5012 37289 5015
rect 4672 4984 37289 5012
rect 4672 4972 4678 4984
rect 37277 4981 37289 4984
rect 37323 4981 37335 5015
rect 38010 5012 38016 5024
rect 37971 4984 38016 5012
rect 37277 4975 37335 4981
rect 38010 4972 38016 4984
rect 38068 4972 38074 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 3234 4604 3240 4616
rect 3195 4576 3240 4604
rect 3234 4564 3240 4576
rect 3292 4604 3298 4616
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3292 4576 3801 4604
rect 3292 4564 3298 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 2774 4264 2780 4276
rect 2735 4236 2780 4264
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 1664 4199 1722 4205
rect 1664 4165 1676 4199
rect 1710 4196 1722 4199
rect 2130 4196 2136 4208
rect 1710 4168 2136 4196
rect 1710 4165 1722 4168
rect 1664 4159 1722 4165
rect 2130 4156 2136 4168
rect 2188 4156 2194 4208
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 37921 4131 37979 4137
rect 37921 4128 37933 4131
rect 37384 4100 37933 4128
rect 37384 3936 37412 4100
rect 37921 4097 37933 4100
rect 37967 4097 37979 4131
rect 37921 4091 37979 4097
rect 38102 3992 38108 4004
rect 38063 3964 38108 3992
rect 38102 3952 38108 3964
rect 38160 3952 38166 4004
rect 37366 3924 37372 3936
rect 37327 3896 37372 3924
rect 37366 3884 37372 3896
rect 37424 3884 37430 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2038 3516 2044 3528
rect 1999 3488 2044 3516
rect 2038 3476 2044 3488
rect 2096 3476 2102 3528
rect 38102 3516 38108 3528
rect 38063 3488 38108 3516
rect 38102 3476 38108 3488
rect 38160 3476 38166 3528
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3380 1915 3383
rect 37366 3380 37372 3392
rect 1903 3352 37372 3380
rect 1903 3349 1915 3352
rect 1857 3343 1915 3349
rect 37366 3340 37372 3352
rect 37424 3340 37430 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 3881 3179 3939 3185
rect 3881 3176 3893 3179
rect 2096 3148 3893 3176
rect 2096 3136 2102 3148
rect 3881 3145 3893 3148
rect 3927 3145 3939 3179
rect 3881 3139 3939 3145
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 2593 3111 2651 3117
rect 2593 3108 2605 3111
rect 2004 3080 2605 3108
rect 2004 3068 2010 3080
rect 2593 3077 2605 3080
rect 2639 3077 2651 3111
rect 2593 3071 2651 3077
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 37372 36728 37424 36780
rect 38016 36635 38068 36644
rect 38016 36601 38025 36635
rect 38025 36601 38059 36635
rect 38059 36601 38068 36635
rect 38016 36592 38068 36601
rect 37372 36567 37424 36576
rect 37372 36533 37381 36567
rect 37381 36533 37415 36567
rect 37415 36533 37424 36567
rect 37372 36524 37424 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 38200 36116 38252 36168
rect 1400 36023 1452 36032
rect 1400 35989 1409 36023
rect 1409 35989 1443 36023
rect 1443 35989 1452 36023
rect 1400 35980 1452 35989
rect 38016 36023 38068 36032
rect 38016 35989 38025 36023
rect 38025 35989 38059 36023
rect 38059 35989 38068 36023
rect 38016 35980 38068 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1400 35683 1452 35692
rect 1400 35649 1409 35683
rect 1409 35649 1443 35683
rect 1443 35649 1452 35683
rect 1400 35640 1452 35649
rect 37740 35640 37792 35692
rect 1492 35504 1544 35556
rect 2504 35436 2556 35488
rect 38016 35479 38068 35488
rect 38016 35445 38025 35479
rect 38025 35445 38059 35479
rect 38059 35445 38068 35479
rect 38016 35436 38068 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1492 35028 1544 35080
rect 38108 35028 38160 35080
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 2044 34935 2096 34944
rect 2044 34901 2053 34935
rect 2053 34901 2087 34935
rect 2087 34901 2096 34935
rect 2044 34892 2096 34901
rect 38016 34935 38068 34944
rect 38016 34901 38025 34935
rect 38025 34901 38059 34935
rect 38059 34901 38068 34935
rect 38016 34892 38068 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1584 34688 1636 34740
rect 19248 34688 19300 34740
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 2044 34552 2096 34604
rect 2228 34595 2280 34604
rect 2228 34561 2237 34595
rect 2237 34561 2271 34595
rect 2271 34561 2280 34595
rect 2228 34552 2280 34561
rect 1676 34348 1728 34400
rect 2044 34391 2096 34400
rect 2044 34357 2053 34391
rect 2053 34357 2087 34391
rect 2087 34357 2096 34391
rect 2044 34348 2096 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 1584 33847 1636 33856
rect 1584 33813 1593 33847
rect 1593 33813 1627 33847
rect 1627 33813 1636 33847
rect 1584 33804 1636 33813
rect 1768 33804 1820 33856
rect 37280 33847 37332 33856
rect 37280 33813 37289 33847
rect 37289 33813 37323 33847
rect 37323 33813 37332 33847
rect 37280 33804 37332 33813
rect 38016 33847 38068 33856
rect 38016 33813 38025 33847
rect 38025 33813 38059 33847
rect 38059 33813 38068 33847
rect 38016 33804 38068 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1584 33600 1636 33652
rect 19156 33600 19208 33652
rect 1584 33464 1636 33516
rect 37464 33464 37516 33516
rect 19984 33328 20036 33380
rect 2872 33260 2924 33312
rect 37464 33260 37516 33312
rect 38016 33303 38068 33312
rect 38016 33269 38025 33303
rect 38025 33269 38059 33303
rect 38059 33269 38068 33303
rect 38016 33260 38068 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2044 33056 2096 33108
rect 1676 32895 1728 32904
rect 1676 32861 1685 32895
rect 1685 32861 1719 32895
rect 1719 32861 1728 32895
rect 1676 32852 1728 32861
rect 2044 32895 2096 32904
rect 2044 32861 2053 32895
rect 2053 32861 2087 32895
rect 2087 32861 2096 32895
rect 2044 32852 2096 32861
rect 2872 32895 2924 32904
rect 2872 32861 2881 32895
rect 2881 32861 2915 32895
rect 2915 32861 2924 32895
rect 2872 32852 2924 32861
rect 1492 32759 1544 32768
rect 1492 32725 1501 32759
rect 1501 32725 1535 32759
rect 1535 32725 1544 32759
rect 1492 32716 1544 32725
rect 37556 32716 37608 32768
rect 38016 32759 38068 32768
rect 38016 32725 38025 32759
rect 38025 32725 38059 32759
rect 38059 32725 38068 32759
rect 38016 32716 38068 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 2044 32512 2096 32564
rect 1768 32444 1820 32496
rect 1492 32376 1544 32428
rect 2136 32376 2188 32428
rect 3056 32419 3108 32428
rect 1860 32308 1912 32360
rect 3056 32385 3065 32419
rect 3065 32385 3099 32419
rect 3099 32385 3108 32419
rect 3056 32376 3108 32385
rect 38292 32376 38344 32428
rect 37372 32240 37424 32292
rect 1676 32172 1728 32224
rect 38016 32215 38068 32224
rect 38016 32181 38025 32215
rect 38025 32181 38059 32215
rect 38059 32181 38068 32215
rect 38016 32172 38068 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2688 31900 2740 31952
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 1492 31696 1544 31748
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1492 31288 1544 31340
rect 2228 31331 2280 31340
rect 2228 31297 2237 31331
rect 2237 31297 2271 31331
rect 2271 31297 2280 31331
rect 2228 31288 2280 31297
rect 37924 31288 37976 31340
rect 38016 31195 38068 31204
rect 38016 31161 38025 31195
rect 38025 31161 38059 31195
rect 38059 31161 38068 31195
rect 38016 31152 38068 31161
rect 1860 31084 1912 31136
rect 2044 31127 2096 31136
rect 2044 31093 2053 31127
rect 2053 31093 2087 31127
rect 2087 31093 2096 31127
rect 2044 31084 2096 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1952 30923 2004 30932
rect 1952 30889 1961 30923
rect 1961 30889 1995 30923
rect 1995 30889 2004 30923
rect 1952 30880 2004 30889
rect 2044 30787 2096 30796
rect 2044 30753 2053 30787
rect 2053 30753 2087 30787
rect 2087 30753 2096 30787
rect 2044 30744 2096 30753
rect 1860 30719 1912 30728
rect 1860 30685 1869 30719
rect 1869 30685 1903 30719
rect 1903 30685 1912 30719
rect 1860 30676 1912 30685
rect 2136 30719 2188 30728
rect 2136 30685 2145 30719
rect 2145 30685 2179 30719
rect 2179 30685 2188 30719
rect 2136 30676 2188 30685
rect 2504 30676 2556 30728
rect 1584 30608 1636 30660
rect 2136 30540 2188 30592
rect 34520 30608 34572 30660
rect 37648 30540 37700 30592
rect 38016 30583 38068 30592
rect 38016 30549 38025 30583
rect 38025 30549 38059 30583
rect 38059 30549 38068 30583
rect 38016 30540 38068 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 34520 30268 34572 30320
rect 1492 30200 1544 30252
rect 2044 30243 2096 30252
rect 2044 30209 2053 30243
rect 2053 30209 2087 30243
rect 2087 30209 2096 30243
rect 2044 30200 2096 30209
rect 2412 30064 2464 30116
rect 2228 30039 2280 30048
rect 2228 30005 2237 30039
rect 2237 30005 2271 30039
rect 2271 30005 2280 30039
rect 2228 29996 2280 30005
rect 38016 30039 38068 30048
rect 38016 30005 38025 30039
rect 38025 30005 38059 30039
rect 38059 30005 38068 30039
rect 38016 29996 38068 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1952 29792 2004 29844
rect 2228 29792 2280 29844
rect 12440 29792 12492 29844
rect 2228 29631 2280 29640
rect 1308 29520 1360 29572
rect 2228 29597 2237 29631
rect 2237 29597 2271 29631
rect 2271 29597 2280 29631
rect 2228 29588 2280 29597
rect 19248 29588 19300 29640
rect 1768 29452 1820 29504
rect 38016 29495 38068 29504
rect 38016 29461 38025 29495
rect 38025 29461 38059 29495
rect 38059 29461 38068 29495
rect 38016 29452 38068 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 2504 29248 2556 29300
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 19156 29112 19208 29164
rect 1584 29044 1636 29096
rect 37280 28976 37332 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 37280 28747 37332 28756
rect 37280 28713 37289 28747
rect 37289 28713 37323 28747
rect 37323 28713 37332 28747
rect 37280 28704 37332 28713
rect 1584 28500 1636 28552
rect 19984 28543 20036 28552
rect 19984 28509 19993 28543
rect 19993 28509 20027 28543
rect 20027 28509 20036 28543
rect 19984 28500 20036 28509
rect 37280 28500 37332 28552
rect 1492 28432 1544 28484
rect 2596 28364 2648 28416
rect 37188 28432 37240 28484
rect 38016 28407 38068 28416
rect 38016 28373 38025 28407
rect 38025 28373 38059 28407
rect 38059 28373 38068 28407
rect 38016 28364 38068 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 37188 28160 37240 28212
rect 1676 28092 1728 28144
rect 1492 28024 1544 28076
rect 2228 28067 2280 28076
rect 2228 28033 2237 28067
rect 2237 28033 2271 28067
rect 2271 28033 2280 28067
rect 2228 28024 2280 28033
rect 37280 27956 37332 28008
rect 1952 27820 2004 27872
rect 2044 27863 2096 27872
rect 2044 27829 2053 27863
rect 2053 27829 2087 27863
rect 2087 27829 2096 27863
rect 38016 27863 38068 27872
rect 2044 27820 2096 27829
rect 38016 27829 38025 27863
rect 38025 27829 38059 27863
rect 38059 27829 38068 27863
rect 38016 27820 38068 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 37280 27591 37332 27600
rect 37280 27557 37289 27591
rect 37289 27557 37323 27591
rect 37323 27557 37332 27591
rect 37280 27548 37332 27557
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 1676 27276 1728 27328
rect 19432 27276 19484 27328
rect 38016 27319 38068 27328
rect 38016 27285 38025 27319
rect 38025 27285 38059 27319
rect 38059 27285 38068 27319
rect 38016 27276 38068 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 2044 27004 2096 27056
rect 1952 26979 2004 26988
rect 1952 26945 1961 26979
rect 1961 26945 1995 26979
rect 1995 26945 2004 26979
rect 1952 26936 2004 26945
rect 1768 26911 1820 26920
rect 1768 26877 1777 26911
rect 1777 26877 1811 26911
rect 1811 26877 1820 26911
rect 1768 26868 1820 26877
rect 2688 26868 2740 26920
rect 1952 26775 2004 26784
rect 1952 26741 1961 26775
rect 1961 26741 1995 26775
rect 1995 26741 2004 26775
rect 1952 26732 2004 26741
rect 2136 26775 2188 26784
rect 2136 26741 2145 26775
rect 2145 26741 2179 26775
rect 2179 26741 2188 26775
rect 2136 26732 2188 26741
rect 2780 26732 2832 26784
rect 38016 26775 38068 26784
rect 38016 26741 38025 26775
rect 38025 26741 38059 26775
rect 38059 26741 38068 26775
rect 38016 26732 38068 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 1952 26528 2004 26580
rect 1768 26460 1820 26512
rect 2596 26392 2648 26444
rect 1492 26324 1544 26376
rect 1676 26324 1728 26376
rect 2044 26367 2096 26376
rect 2044 26333 2053 26367
rect 2053 26333 2087 26367
rect 2087 26333 2096 26367
rect 2044 26324 2096 26333
rect 2780 26324 2832 26376
rect 12440 26324 12492 26376
rect 16580 26256 16632 26308
rect 37188 26256 37240 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2596 26027 2648 26036
rect 2596 25993 2605 26027
rect 2605 25993 2639 26027
rect 2639 25993 2648 26027
rect 2596 25984 2648 25993
rect 37188 25984 37240 26036
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 2412 25712 2464 25764
rect 37188 25712 37240 25764
rect 38016 25755 38068 25764
rect 38016 25721 38025 25755
rect 38025 25721 38059 25755
rect 38059 25721 38068 25755
rect 38016 25712 38068 25721
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 1952 25644 2004 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1584 25440 1636 25492
rect 13820 25440 13872 25492
rect 37188 25440 37240 25492
rect 1492 25236 1544 25288
rect 2504 25168 2556 25220
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 2136 25143 2188 25152
rect 2136 25109 2145 25143
rect 2145 25109 2179 25143
rect 2179 25109 2188 25143
rect 2136 25100 2188 25109
rect 33140 25168 33192 25220
rect 38016 25143 38068 25152
rect 38016 25109 38025 25143
rect 38025 25109 38059 25143
rect 38059 25109 38068 25143
rect 38016 25100 38068 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1584 24896 1636 24948
rect 19984 24896 20036 24948
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 1952 24760 2004 24812
rect 2136 24760 2188 24812
rect 33140 24760 33192 24812
rect 1676 24556 1728 24608
rect 2780 24599 2832 24608
rect 2780 24565 2789 24599
rect 2789 24565 2823 24599
rect 2823 24565 2832 24599
rect 2780 24556 2832 24565
rect 17776 24556 17828 24608
rect 38016 24599 38068 24608
rect 38016 24565 38025 24599
rect 38025 24565 38059 24599
rect 38059 24565 38068 24599
rect 38016 24556 38068 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1584 24352 1636 24404
rect 1768 24259 1820 24268
rect 1768 24225 1777 24259
rect 1777 24225 1811 24259
rect 1811 24225 1820 24259
rect 1768 24216 1820 24225
rect 1676 24191 1728 24200
rect 1676 24157 1685 24191
rect 1685 24157 1719 24191
rect 1719 24157 1728 24191
rect 1676 24148 1728 24157
rect 2780 24191 2832 24200
rect 2412 24012 2464 24064
rect 2780 24157 2789 24191
rect 2789 24157 2823 24191
rect 2823 24157 2832 24191
rect 2780 24148 2832 24157
rect 19800 24191 19852 24200
rect 19800 24157 19809 24191
rect 19809 24157 19843 24191
rect 19843 24157 19852 24191
rect 19800 24148 19852 24157
rect 38016 24055 38068 24064
rect 38016 24021 38025 24055
rect 38025 24021 38059 24055
rect 38059 24021 38068 24055
rect 38016 24012 38068 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 2228 23783 2280 23792
rect 2228 23749 2237 23783
rect 2237 23749 2271 23783
rect 2271 23749 2280 23783
rect 2228 23740 2280 23749
rect 1492 23672 1544 23724
rect 2412 23715 2464 23724
rect 2412 23681 2421 23715
rect 2421 23681 2455 23715
rect 2455 23681 2464 23715
rect 2412 23672 2464 23681
rect 2504 23715 2556 23724
rect 2504 23681 2513 23715
rect 2513 23681 2547 23715
rect 2547 23681 2556 23715
rect 2504 23672 2556 23681
rect 19432 23672 19484 23724
rect 2044 23468 2096 23520
rect 4620 23468 4672 23520
rect 37280 23468 37332 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 37280 23307 37332 23316
rect 37280 23273 37289 23307
rect 37289 23273 37323 23307
rect 37323 23273 37332 23307
rect 37280 23264 37332 23273
rect 1492 23196 1544 23248
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 4620 23060 4672 23112
rect 16580 23060 16632 23112
rect 37280 23060 37332 23112
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 4620 22924 4672 22976
rect 31024 22992 31076 23044
rect 38016 22967 38068 22976
rect 38016 22933 38025 22967
rect 38025 22933 38059 22967
rect 38059 22933 38068 22967
rect 38016 22924 38068 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1584 22720 1636 22772
rect 17868 22720 17920 22772
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 13820 22584 13872 22636
rect 31024 22584 31076 22636
rect 1768 22380 1820 22432
rect 37280 22380 37332 22432
rect 38016 22423 38068 22432
rect 38016 22389 38025 22423
rect 38025 22389 38059 22423
rect 38059 22389 38068 22423
rect 38016 22380 38068 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 37280 22083 37332 22092
rect 37280 22049 37289 22083
rect 37289 22049 37323 22083
rect 37323 22049 37332 22083
rect 37280 22040 37332 22049
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 17960 21836 18012 21888
rect 38016 21879 38068 21888
rect 38016 21845 38025 21879
rect 38025 21845 38059 21879
rect 38059 21845 38068 21879
rect 38016 21836 38068 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 19984 21539 20036 21548
rect 19984 21505 19993 21539
rect 19993 21505 20027 21539
rect 20027 21505 20036 21539
rect 19984 21496 20036 21505
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 2780 21292 2832 21344
rect 38016 21335 38068 21344
rect 38016 21301 38025 21335
rect 38025 21301 38059 21335
rect 38059 21301 38068 21335
rect 38016 21292 38068 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1492 20952 1544 21004
rect 2780 20952 2832 21004
rect 2228 20927 2280 20936
rect 2228 20893 2237 20927
rect 2237 20893 2271 20927
rect 2271 20893 2280 20927
rect 2228 20884 2280 20893
rect 17776 20884 17828 20936
rect 18972 20816 19024 20868
rect 1952 20748 2004 20800
rect 19432 20791 19484 20800
rect 19432 20757 19441 20791
rect 19441 20757 19475 20791
rect 19475 20757 19484 20791
rect 19432 20748 19484 20757
rect 33140 20816 33192 20868
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 33140 20544 33192 20596
rect 1584 20476 1636 20528
rect 17868 20476 17920 20528
rect 1952 20451 2004 20460
rect 1952 20417 1961 20451
rect 1961 20417 1995 20451
rect 1995 20417 2004 20451
rect 1952 20408 2004 20417
rect 2872 20408 2924 20460
rect 18972 20451 19024 20460
rect 18972 20417 18981 20451
rect 18981 20417 19015 20451
rect 19015 20417 19024 20451
rect 18972 20408 19024 20417
rect 19432 20408 19484 20460
rect 1768 20383 1820 20392
rect 1768 20349 1777 20383
rect 1777 20349 1811 20383
rect 1811 20349 1820 20383
rect 1768 20340 1820 20349
rect 19892 20315 19944 20324
rect 19892 20281 19901 20315
rect 19901 20281 19935 20315
rect 19935 20281 19944 20315
rect 19892 20272 19944 20281
rect 31024 20272 31076 20324
rect 38016 20315 38068 20324
rect 38016 20281 38025 20315
rect 38025 20281 38059 20315
rect 38059 20281 38068 20315
rect 38016 20272 38068 20281
rect 1584 20204 1636 20256
rect 2044 20204 2096 20256
rect 2780 20247 2832 20256
rect 2780 20213 2789 20247
rect 2789 20213 2823 20247
rect 2823 20213 2832 20247
rect 2780 20204 2832 20213
rect 19156 20247 19208 20256
rect 19156 20213 19165 20247
rect 19165 20213 19199 20247
rect 19199 20213 19208 20247
rect 19156 20204 19208 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 2504 20000 2556 20052
rect 19156 20000 19208 20052
rect 31760 20000 31812 20052
rect 2780 19932 2832 19984
rect 21088 19932 21140 19984
rect 1768 19864 1820 19916
rect 2044 19796 2096 19848
rect 2228 19796 2280 19848
rect 2780 19839 2832 19848
rect 2780 19805 2789 19839
rect 2789 19805 2823 19839
rect 2823 19805 2832 19839
rect 2780 19796 2832 19805
rect 18512 19796 18564 19848
rect 14464 19728 14516 19780
rect 17868 19660 17920 19712
rect 18512 19660 18564 19712
rect 20628 19771 20680 19780
rect 20628 19737 20637 19771
rect 20637 19737 20671 19771
rect 20671 19737 20680 19771
rect 20628 19728 20680 19737
rect 31024 19796 31076 19848
rect 37648 19660 37700 19712
rect 38016 19703 38068 19712
rect 38016 19669 38025 19703
rect 38025 19669 38059 19703
rect 38059 19669 38068 19703
rect 38016 19660 38068 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 2228 19499 2280 19508
rect 2228 19465 2237 19499
rect 2237 19465 2271 19499
rect 2271 19465 2280 19499
rect 2228 19456 2280 19465
rect 17960 19499 18012 19508
rect 17960 19465 17969 19499
rect 17969 19465 18003 19499
rect 18003 19465 18012 19499
rect 17960 19456 18012 19465
rect 2780 19431 2832 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2044 19363 2096 19372
rect 2044 19329 2053 19363
rect 2053 19329 2087 19363
rect 2087 19329 2096 19363
rect 2044 19320 2096 19329
rect 2780 19397 2789 19431
rect 2789 19397 2823 19431
rect 2823 19397 2832 19431
rect 2780 19388 2832 19397
rect 27528 19456 27580 19508
rect 20352 19320 20404 19372
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 18420 19159 18472 19168
rect 18420 19125 18429 19159
rect 18429 19125 18463 19159
rect 18463 19125 18472 19159
rect 18420 19116 18472 19125
rect 38292 19184 38344 19236
rect 37464 19116 37516 19168
rect 38016 19159 38068 19168
rect 38016 19125 38025 19159
rect 38025 19125 38059 19159
rect 38059 19125 38068 19159
rect 38016 19116 38068 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1860 18955 1912 18964
rect 1860 18921 1869 18955
rect 1869 18921 1903 18955
rect 1903 18921 1912 18955
rect 1860 18912 1912 18921
rect 2044 18912 2096 18964
rect 21088 18912 21140 18964
rect 31760 18912 31812 18964
rect 1952 18751 2004 18760
rect 1952 18717 1961 18751
rect 1961 18717 1995 18751
rect 1995 18717 2004 18751
rect 1952 18708 2004 18717
rect 20076 18708 20128 18760
rect 2320 18640 2372 18692
rect 20352 18615 20404 18624
rect 20352 18581 20361 18615
rect 20361 18581 20395 18615
rect 20395 18581 20404 18615
rect 20352 18572 20404 18581
rect 37372 18572 37424 18624
rect 38016 18615 38068 18624
rect 38016 18581 38025 18615
rect 38025 18581 38059 18615
rect 38059 18581 38068 18615
rect 38016 18572 38068 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 17960 18096 18012 18148
rect 20720 18096 20772 18148
rect 20076 18028 20128 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1952 17824 2004 17876
rect 1400 17756 1452 17808
rect 1492 17620 1544 17672
rect 17868 17620 17920 17672
rect 27528 17620 27580 17672
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 38200 17552 38252 17604
rect 31024 17484 31076 17536
rect 38016 17527 38068 17536
rect 38016 17493 38025 17527
rect 38025 17493 38059 17527
rect 38059 17493 38068 17527
rect 38016 17484 38068 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1492 17280 1544 17332
rect 13912 17212 13964 17264
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 18604 17008 18656 17060
rect 15108 16940 15160 16992
rect 31024 17144 31076 17196
rect 38108 17008 38160 17060
rect 37740 16940 37792 16992
rect 38016 16983 38068 16992
rect 38016 16949 38025 16983
rect 38025 16949 38059 16983
rect 38059 16949 38068 16983
rect 38016 16940 38068 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 20720 16779 20772 16788
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 1492 16532 1544 16584
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 17960 16532 18012 16584
rect 19248 16532 19300 16584
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 2228 16439 2280 16448
rect 2228 16405 2237 16439
rect 2237 16405 2271 16439
rect 2271 16405 2280 16439
rect 2228 16396 2280 16405
rect 37188 16396 37240 16448
rect 38016 16439 38068 16448
rect 38016 16405 38025 16439
rect 38025 16405 38059 16439
rect 38059 16405 38068 16439
rect 38016 16396 38068 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 1584 16192 1636 16244
rect 1492 16124 1544 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 19248 16192 19300 16244
rect 37188 16192 37240 16244
rect 15108 15920 15160 15972
rect 33140 15920 33192 15972
rect 38016 15895 38068 15904
rect 38016 15861 38025 15895
rect 38025 15861 38059 15895
rect 38059 15861 38068 15895
rect 38016 15852 38068 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1492 15648 1544 15700
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 13912 15376 13964 15428
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 33140 15104 33192 15156
rect 2228 15036 2280 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 19984 14832 20036 14884
rect 37280 14900 37332 14952
rect 38016 14875 38068 14884
rect 38016 14841 38025 14875
rect 38025 14841 38059 14875
rect 38059 14841 38068 14875
rect 38016 14832 38068 14841
rect 19432 14764 19484 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1492 14560 1544 14612
rect 37280 14603 37332 14612
rect 37280 14569 37289 14603
rect 37289 14569 37323 14603
rect 37323 14569 37332 14603
rect 37280 14560 37332 14569
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 19984 14399 20036 14408
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 37188 14220 37240 14272
rect 38016 14263 38068 14272
rect 38016 14229 38025 14263
rect 38025 14229 38059 14263
rect 38059 14229 38068 14263
rect 38016 14220 38068 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 37188 14016 37240 14068
rect 20352 13948 20404 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 19432 13880 19484 13932
rect 37188 13812 37240 13864
rect 2228 13719 2280 13728
rect 2228 13685 2237 13719
rect 2237 13685 2271 13719
rect 2271 13685 2280 13719
rect 2228 13676 2280 13685
rect 38016 13719 38068 13728
rect 38016 13685 38025 13719
rect 38025 13685 38059 13719
rect 38059 13685 38068 13719
rect 38016 13676 38068 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 37188 13472 37240 13524
rect 19340 13336 19392 13388
rect 2136 13268 2188 13320
rect 2780 13268 2832 13320
rect 15200 13132 15252 13184
rect 38016 13175 38068 13184
rect 38016 13141 38025 13175
rect 38025 13141 38059 13175
rect 38059 13141 38068 13175
rect 38016 13132 38068 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 2228 12928 2280 12980
rect 2780 12903 2832 12912
rect 2780 12869 2789 12903
rect 2789 12869 2823 12903
rect 2823 12869 2832 12903
rect 2780 12860 2832 12869
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 18420 12724 18472 12776
rect 37004 12588 37056 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2136 12427 2188 12436
rect 2136 12393 2145 12427
rect 2145 12393 2179 12427
rect 2179 12393 2188 12427
rect 2136 12384 2188 12393
rect 2228 12384 2280 12436
rect 37004 12384 37056 12436
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 15200 12180 15252 12232
rect 15292 12112 15344 12164
rect 37188 12044 37240 12096
rect 38016 12087 38068 12096
rect 38016 12053 38025 12087
rect 38025 12053 38059 12087
rect 38059 12053 38068 12087
rect 38016 12044 38068 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 37188 11840 37240 11892
rect 14464 11704 14516 11756
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 38016 11543 38068 11552
rect 38016 11509 38025 11543
rect 38025 11509 38059 11543
rect 38059 11509 38068 11543
rect 38016 11500 38068 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1492 11296 1544 11348
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 38016 11271 38068 11280
rect 38016 11237 38025 11271
rect 38025 11237 38059 11271
rect 38059 11237 38068 11271
rect 38016 11228 38068 11237
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 19708 10480 19760 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 37280 10455 37332 10464
rect 37280 10421 37289 10455
rect 37289 10421 37323 10455
rect 37323 10421 37332 10455
rect 37280 10412 37332 10421
rect 38016 10455 38068 10464
rect 38016 10421 38025 10455
rect 38025 10421 38059 10455
rect 38059 10421 38068 10455
rect 38016 10412 38068 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1584 10208 1636 10260
rect 13820 10208 13872 10260
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 18512 10004 18564 10056
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 37280 9868 37332 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 1400 9664 1452 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 19708 9571 19760 9580
rect 19708 9537 19717 9571
rect 19717 9537 19751 9571
rect 19751 9537 19760 9571
rect 19708 9528 19760 9537
rect 38016 9435 38068 9444
rect 38016 9401 38025 9435
rect 38025 9401 38059 9435
rect 38059 9401 38068 9435
rect 38016 9392 38068 9401
rect 18420 9324 18472 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1492 9120 1544 9172
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 19708 8916 19760 8968
rect 13820 8848 13872 8900
rect 20628 8848 20680 8900
rect 19432 8780 19484 8832
rect 37280 8823 37332 8832
rect 37280 8789 37289 8823
rect 37289 8789 37323 8823
rect 37323 8789 37332 8823
rect 37280 8780 37332 8789
rect 38016 8823 38068 8832
rect 38016 8789 38025 8823
rect 38025 8789 38059 8823
rect 38059 8789 38068 8823
rect 38016 8780 38068 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 15292 8576 15344 8628
rect 2320 8551 2372 8560
rect 2320 8517 2329 8551
rect 2329 8517 2363 8551
rect 2363 8517 2372 8551
rect 2320 8508 2372 8517
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 18604 8372 18656 8424
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 19432 8372 19484 8424
rect 37280 8508 37332 8560
rect 37372 8440 37424 8492
rect 38016 8347 38068 8356
rect 38016 8313 38025 8347
rect 38025 8313 38059 8347
rect 38059 8313 38068 8347
rect 38016 8304 38068 8313
rect 20628 8236 20680 8288
rect 21272 8236 21324 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1400 8032 1452 8084
rect 18420 8032 18472 8084
rect 2320 7964 2372 8016
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 19432 7828 19484 7880
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 20628 7692 20680 7744
rect 37372 7760 37424 7812
rect 38016 7735 38068 7744
rect 38016 7701 38025 7735
rect 38025 7701 38059 7735
rect 38059 7701 38068 7735
rect 38016 7692 38068 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 18604 7531 18656 7540
rect 18604 7497 18613 7531
rect 18613 7497 18647 7531
rect 18647 7497 18656 7531
rect 18604 7488 18656 7497
rect 1768 7352 1820 7404
rect 19432 7352 19484 7404
rect 20076 7352 20128 7404
rect 20628 7395 20680 7404
rect 20628 7361 20637 7395
rect 20637 7361 20671 7395
rect 20671 7361 20680 7395
rect 20628 7352 20680 7361
rect 19524 7191 19576 7200
rect 19524 7157 19533 7191
rect 19533 7157 19567 7191
rect 19567 7157 19576 7191
rect 19524 7148 19576 7157
rect 37832 7148 37884 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 2780 6740 2832 6792
rect 19524 6740 19576 6792
rect 37832 6783 37884 6792
rect 37832 6749 37841 6783
rect 37841 6749 37875 6783
rect 37875 6749 37884 6783
rect 37832 6740 37884 6749
rect 37832 6604 37884 6656
rect 38016 6647 38068 6656
rect 38016 6613 38025 6647
rect 38025 6613 38059 6647
rect 38059 6613 38068 6647
rect 38016 6604 38068 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2136 6264 2188 6316
rect 20076 6264 20128 6316
rect 37832 6307 37884 6316
rect 37832 6273 37841 6307
rect 37841 6273 37875 6307
rect 37875 6273 37884 6307
rect 37832 6264 37884 6273
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 37832 6060 37884 6112
rect 38016 6103 38068 6112
rect 38016 6069 38025 6103
rect 38025 6069 38059 6103
rect 38059 6069 38068 6103
rect 38016 6060 38068 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 37832 5695 37884 5704
rect 37832 5661 37841 5695
rect 37841 5661 37875 5695
rect 37875 5661 37884 5695
rect 37832 5652 37884 5661
rect 1400 5584 1452 5636
rect 1952 5584 2004 5636
rect 38016 5559 38068 5568
rect 38016 5525 38025 5559
rect 38025 5525 38059 5559
rect 38059 5525 38068 5559
rect 38016 5516 38068 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1768 5312 1820 5364
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 1308 5176 1360 5228
rect 1860 5176 1912 5228
rect 2780 5176 2832 5228
rect 4620 4972 4672 5024
rect 38016 5015 38068 5024
rect 38016 4981 38025 5015
rect 38025 4981 38059 5015
rect 38059 4981 38068 5015
rect 38016 4972 38068 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 2780 4224 2832 4233
rect 2136 4156 2188 4208
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 38108 3995 38160 4004
rect 38108 3961 38117 3995
rect 38117 3961 38151 3995
rect 38151 3961 38160 3995
rect 38108 3952 38160 3961
rect 37372 3927 37424 3936
rect 37372 3893 37381 3927
rect 37381 3893 37415 3927
rect 37415 3893 37424 3927
rect 37372 3884 37424 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 38108 3519 38160 3528
rect 38108 3485 38117 3519
rect 38117 3485 38151 3519
rect 38151 3485 38160 3519
rect 38108 3476 38160 3485
rect 37372 3340 37424 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2044 3136 2096 3188
rect 1952 3068 2004 3120
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 37372 36780 37424 36786
rect 37372 36722 37424 36728
rect 37384 36582 37412 36722
rect 38014 36680 38070 36689
rect 38014 36615 38016 36624
rect 38068 36615 38070 36624
rect 38016 36586 38068 36592
rect 37372 36576 37424 36582
rect 37372 36518 37424 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 1400 36032 1452 36038
rect 1400 35974 1452 35980
rect 1412 35698 1440 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 1412 34921 1440 35634
rect 1492 35556 1544 35562
rect 1492 35498 1544 35504
rect 1504 35086 1532 35498
rect 2504 35488 2556 35494
rect 2504 35430 2556 35436
rect 1492 35080 1544 35086
rect 1492 35022 1544 35028
rect 1398 34912 1454 34921
rect 1398 34847 1454 34856
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1412 34490 1440 34546
rect 1320 34462 1440 34490
rect 1320 33697 1348 34462
rect 1504 34105 1532 35022
rect 1584 34944 1636 34950
rect 1584 34886 1636 34892
rect 2044 34944 2096 34950
rect 2044 34886 2096 34892
rect 1596 34746 1624 34886
rect 1584 34740 1636 34746
rect 1584 34682 1636 34688
rect 2056 34610 2084 34886
rect 2044 34604 2096 34610
rect 2044 34546 2096 34552
rect 2228 34604 2280 34610
rect 2228 34546 2280 34552
rect 2240 34513 2268 34546
rect 2226 34504 2282 34513
rect 2226 34439 2282 34448
rect 1676 34400 1728 34406
rect 1676 34342 1728 34348
rect 2044 34400 2096 34406
rect 2044 34342 2096 34348
rect 1490 34096 1546 34105
rect 1490 34031 1546 34040
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1306 33688 1362 33697
rect 1306 33623 1362 33632
rect 1412 33289 1440 33934
rect 1584 33856 1636 33862
rect 1584 33798 1636 33804
rect 1596 33658 1624 33798
rect 1584 33652 1636 33658
rect 1584 33594 1636 33600
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1398 33280 1454 33289
rect 1398 33215 1454 33224
rect 1492 32768 1544 32774
rect 1492 32710 1544 32716
rect 1504 32434 1532 32710
rect 1596 32473 1624 33458
rect 1688 32910 1716 34342
rect 1768 33856 1820 33862
rect 1768 33798 1820 33804
rect 1676 32904 1728 32910
rect 1676 32846 1728 32852
rect 1780 32502 1808 33798
rect 2056 33114 2084 34342
rect 2044 33108 2096 33114
rect 2044 33050 2096 33056
rect 2044 32904 2096 32910
rect 2044 32846 2096 32852
rect 2056 32570 2084 32846
rect 2044 32564 2096 32570
rect 2044 32506 2096 32512
rect 1768 32496 1820 32502
rect 1582 32464 1638 32473
rect 1492 32428 1544 32434
rect 1768 32438 1820 32444
rect 1582 32399 1638 32408
rect 1492 32370 1544 32376
rect 1676 32224 1728 32230
rect 1676 32166 1728 32172
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 30841 1440 31758
rect 1492 31748 1544 31754
rect 1492 31690 1544 31696
rect 1504 31346 1532 31690
rect 1492 31340 1544 31346
rect 1492 31282 1544 31288
rect 1398 30832 1454 30841
rect 1398 30767 1454 30776
rect 1504 30433 1532 31282
rect 1584 30660 1636 30666
rect 1584 30602 1636 30608
rect 1490 30424 1546 30433
rect 1490 30359 1546 30368
rect 1596 30274 1624 30602
rect 1504 30258 1624 30274
rect 1492 30252 1624 30258
rect 1544 30246 1624 30252
rect 1492 30194 1544 30200
rect 1308 29572 1360 29578
rect 1308 29514 1360 29520
rect 1320 28801 1348 29514
rect 1504 29209 1532 30194
rect 1490 29200 1546 29209
rect 1400 29164 1452 29170
rect 1490 29135 1546 29144
rect 1400 29106 1452 29112
rect 1306 28792 1362 28801
rect 1306 28727 1362 28736
rect 1412 28393 1440 29106
rect 1584 29096 1636 29102
rect 1584 29038 1636 29044
rect 1596 28558 1624 29038
rect 1584 28552 1636 28558
rect 1584 28494 1636 28500
rect 1492 28484 1544 28490
rect 1492 28426 1544 28432
rect 1398 28384 1454 28393
rect 1398 28319 1454 28328
rect 1504 28082 1532 28426
rect 1492 28076 1544 28082
rect 1492 28018 1544 28024
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 26761 1440 27406
rect 1504 27169 1532 28018
rect 1596 27577 1624 28494
rect 1688 28150 1716 32166
rect 1780 31657 1808 32438
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 1860 32360 1912 32366
rect 1860 32302 1912 32308
rect 1766 31648 1822 31657
rect 1766 31583 1822 31592
rect 1872 31226 1900 32302
rect 1780 31198 1900 31226
rect 1780 29594 1808 31198
rect 1860 31136 1912 31142
rect 1860 31078 1912 31084
rect 2044 31136 2096 31142
rect 2044 31078 2096 31084
rect 1872 30734 1900 31078
rect 1952 30932 2004 30938
rect 1952 30874 2004 30880
rect 1860 30728 1912 30734
rect 1860 30670 1912 30676
rect 1964 29850 1992 30874
rect 2056 30802 2084 31078
rect 2044 30796 2096 30802
rect 2044 30738 2096 30744
rect 2148 30734 2176 32370
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 2240 31249 2268 31282
rect 2226 31240 2282 31249
rect 2226 31175 2282 31184
rect 2516 30734 2544 35430
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19248 34740 19300 34746
rect 19248 34682 19300 34688
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19156 33652 19208 33658
rect 19156 33594 19208 33600
rect 2872 33312 2924 33318
rect 2872 33254 2924 33260
rect 2884 32910 2912 33254
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 2872 32904 2924 32910
rect 2870 32872 2872 32881
rect 2924 32872 2926 32881
rect 2870 32807 2926 32816
rect 3056 32428 3108 32434
rect 3056 32370 3108 32376
rect 3068 32065 3096 32370
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 3054 32056 3110 32065
rect 4214 32059 4522 32068
rect 3054 31991 3110 32000
rect 2688 31952 2740 31958
rect 2688 31894 2740 31900
rect 2136 30728 2188 30734
rect 2136 30670 2188 30676
rect 2504 30728 2556 30734
rect 2504 30670 2556 30676
rect 2136 30592 2188 30598
rect 2136 30534 2188 30540
rect 2044 30252 2096 30258
rect 2044 30194 2096 30200
rect 2056 30025 2084 30194
rect 2042 30016 2098 30025
rect 2042 29951 2098 29960
rect 1952 29844 2004 29850
rect 1952 29786 2004 29792
rect 1780 29566 1900 29594
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 1676 28144 1728 28150
rect 1676 28086 1728 28092
rect 1582 27568 1638 27577
rect 1582 27503 1638 27512
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1490 27160 1546 27169
rect 1490 27095 1546 27104
rect 1398 26752 1454 26761
rect 1398 26687 1454 26696
rect 1688 26382 1716 27270
rect 1780 26926 1808 29446
rect 1768 26920 1820 26926
rect 1768 26862 1820 26868
rect 1768 26512 1820 26518
rect 1768 26454 1820 26460
rect 1492 26376 1544 26382
rect 1492 26318 1544 26324
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1412 25129 1440 25842
rect 1504 25537 1532 26318
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1490 25528 1546 25537
rect 1596 25498 1624 25638
rect 1490 25463 1546 25472
rect 1584 25492 1636 25498
rect 1584 25434 1636 25440
rect 1492 25288 1544 25294
rect 1492 25230 1544 25236
rect 1398 25120 1454 25129
rect 1398 25055 1454 25064
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1412 23497 1440 24754
rect 1504 24313 1532 25230
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 24954 1624 25094
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1676 24608 1728 24614
rect 1676 24550 1728 24556
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1490 24304 1546 24313
rect 1490 24239 1546 24248
rect 1596 23866 1624 24346
rect 1688 24206 1716 24550
rect 1780 24274 1808 26454
rect 1768 24268 1820 24274
rect 1768 24210 1820 24216
rect 1676 24200 1728 24206
rect 1676 24142 1728 24148
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1398 23488 1454 23497
rect 1398 23423 1454 23432
rect 1504 23254 1532 23666
rect 1492 23248 1544 23254
rect 1492 23190 1544 23196
rect 1400 23112 1452 23118
rect 1504 23089 1532 23190
rect 1400 23054 1452 23060
rect 1490 23080 1546 23089
rect 1412 22817 1440 23054
rect 1490 23015 1546 23024
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1398 22808 1454 22817
rect 1596 22778 1624 22918
rect 1398 22743 1454 22752
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22273 1440 22578
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 1398 22264 1454 22273
rect 1398 22199 1454 22208
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21865 1440 21966
rect 1398 21856 1454 21865
rect 1398 21791 1454 21800
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21457 1440 21490
rect 1398 21448 1454 21457
rect 1398 21383 1454 21392
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1490 21040 1546 21049
rect 1490 20975 1492 20984
rect 1544 20975 1546 20984
rect 1492 20946 1544 20952
rect 1596 20534 1624 21286
rect 1584 20528 1636 20534
rect 1584 20470 1636 20476
rect 1780 20398 1808 22374
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1398 19816 1454 19825
rect 1398 19751 1454 19760
rect 1412 19378 1440 19751
rect 1596 19514 1624 20198
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1398 18592 1454 18601
rect 1398 18527 1454 18536
rect 1412 18290 1440 18527
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17814 1440 18226
rect 1490 18184 1546 18193
rect 1490 18119 1546 18128
rect 1400 17808 1452 17814
rect 1400 17750 1452 17756
rect 1504 17678 1532 18119
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1398 17368 1454 17377
rect 1504 17338 1532 17614
rect 1398 17303 1454 17312
rect 1492 17332 1544 17338
rect 1412 17202 1440 17303
rect 1492 17274 1544 17280
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1398 16960 1454 16969
rect 1398 16895 1454 16904
rect 1412 16574 1440 16895
rect 1492 16584 1544 16590
rect 1412 16546 1492 16574
rect 1780 16574 1808 19858
rect 1872 18970 1900 29566
rect 1952 27872 2004 27878
rect 1952 27814 2004 27820
rect 2044 27872 2096 27878
rect 2044 27814 2096 27820
rect 2148 27826 2176 30534
rect 2412 30116 2464 30122
rect 2412 30058 2464 30064
rect 2228 30048 2280 30054
rect 2228 29990 2280 29996
rect 2240 29850 2268 29990
rect 2228 29844 2280 29850
rect 2228 29786 2280 29792
rect 2228 29640 2280 29646
rect 2226 29608 2228 29617
rect 2280 29608 2282 29617
rect 2226 29543 2282 29552
rect 2228 28076 2280 28082
rect 2228 28018 2280 28024
rect 2240 27985 2268 28018
rect 2226 27976 2282 27985
rect 2226 27911 2282 27920
rect 1964 26994 1992 27814
rect 2056 27062 2084 27814
rect 2148 27798 2268 27826
rect 2044 27056 2096 27062
rect 2044 26998 2096 27004
rect 1952 26988 2004 26994
rect 1952 26930 2004 26936
rect 1952 26784 2004 26790
rect 1952 26726 2004 26732
rect 2136 26784 2188 26790
rect 2136 26726 2188 26732
rect 1964 26586 1992 26726
rect 1952 26580 2004 26586
rect 1952 26522 2004 26528
rect 2044 26376 2096 26382
rect 2044 26318 2096 26324
rect 2056 25945 2084 26318
rect 2042 25936 2098 25945
rect 2042 25871 2098 25880
rect 1952 25696 2004 25702
rect 1952 25638 2004 25644
rect 1964 24818 1992 25638
rect 2148 25242 2176 26726
rect 2056 25214 2176 25242
rect 1952 24812 2004 24818
rect 1952 24754 2004 24760
rect 2056 23526 2084 25214
rect 2136 25152 2188 25158
rect 2136 25094 2188 25100
rect 2148 24818 2176 25094
rect 2136 24812 2188 24818
rect 2136 24754 2188 24760
rect 2148 24721 2176 24754
rect 2134 24712 2190 24721
rect 2134 24647 2190 24656
rect 2240 23798 2268 27798
rect 2424 25770 2452 30058
rect 2504 29300 2556 29306
rect 2504 29242 2556 29248
rect 2412 25764 2464 25770
rect 2412 25706 2464 25712
rect 2516 25226 2544 29242
rect 2596 28416 2648 28422
rect 2596 28358 2648 28364
rect 2608 27713 2636 28358
rect 2594 27704 2650 27713
rect 2594 27639 2650 27648
rect 2700 26926 2728 31894
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 12440 29844 12492 29850
rect 12440 29786 12492 29792
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 2688 26920 2740 26926
rect 2688 26862 2740 26868
rect 2780 26784 2832 26790
rect 2780 26726 2832 26732
rect 2596 26444 2648 26450
rect 2596 26386 2648 26392
rect 2608 26353 2636 26386
rect 2792 26382 2820 26726
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 12452 26382 12480 29786
rect 19168 29170 19196 33594
rect 19260 29646 19288 34682
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 37280 33856 37332 33862
rect 37280 33798 37332 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19984 33380 20036 33386
rect 19984 33322 20036 33328
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19996 28558 20024 33322
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 37292 31362 37320 33798
rect 37384 32298 37412 36518
rect 38200 36168 38252 36174
rect 38200 36110 38252 36116
rect 38016 36032 38068 36038
rect 38014 36000 38016 36009
rect 38068 36000 38070 36009
rect 38014 35935 38070 35944
rect 37740 35692 37792 35698
rect 37740 35634 37792 35640
rect 37464 33516 37516 33522
rect 37464 33458 37516 33464
rect 37476 33318 37504 33458
rect 37464 33312 37516 33318
rect 37464 33254 37516 33260
rect 37372 32292 37424 32298
rect 37372 32234 37424 32240
rect 37292 31334 37412 31362
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34520 30660 34572 30666
rect 34520 30602 34572 30608
rect 34532 30326 34560 30602
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 37280 29028 37332 29034
rect 37280 28970 37332 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 37292 28762 37320 28970
rect 37280 28756 37332 28762
rect 37280 28698 37332 28704
rect 37292 28558 37320 28698
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 37280 28552 37332 28558
rect 37280 28494 37332 28500
rect 37188 28484 37240 28490
rect 37188 28426 37240 28432
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 37200 28218 37228 28426
rect 37188 28212 37240 28218
rect 37188 28154 37240 28160
rect 37280 28008 37332 28014
rect 37280 27950 37332 27956
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 37292 27606 37320 27950
rect 37280 27600 37332 27606
rect 37280 27542 37332 27548
rect 19432 27328 19484 27334
rect 19432 27270 19484 27276
rect 2780 26376 2832 26382
rect 2594 26344 2650 26353
rect 2780 26318 2832 26324
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 2594 26279 2650 26288
rect 16580 26308 16632 26314
rect 2608 26042 2636 26279
rect 16580 26250 16632 26256
rect 2596 26036 2648 26042
rect 2596 25978 2648 25984
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 13820 25492 13872 25498
rect 13820 25434 13872 25440
rect 2504 25220 2556 25226
rect 2504 25162 2556 25168
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2792 24206 2820 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2412 24064 2464 24070
rect 2412 24006 2464 24012
rect 2228 23792 2280 23798
rect 2228 23734 2280 23740
rect 2424 23730 2452 24006
rect 2792 23905 2820 24142
rect 2778 23896 2834 23905
rect 2778 23831 2834 23840
rect 2412 23724 2464 23730
rect 2412 23666 2464 23672
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1964 20466 1992 20742
rect 2240 20641 2268 20878
rect 2226 20632 2282 20641
rect 2226 20567 2282 20576
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1964 18766 1992 19994
rect 2056 19854 2084 20198
rect 2516 20058 2544 23666
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23118 4660 23462
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2792 21010 2820 21286
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2780 20256 2832 20262
rect 2884 20233 2912 20402
rect 2780 20198 2832 20204
rect 2870 20224 2926 20233
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 2792 19990 2820 20198
rect 2870 20159 2926 20168
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 2780 19984 2832 19990
rect 2780 19926 2832 19932
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2240 19514 2268 19790
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 2792 19446 2820 19790
rect 2780 19440 2832 19446
rect 2778 19408 2780 19417
rect 2832 19408 2834 19417
rect 2044 19372 2096 19378
rect 2778 19343 2834 19352
rect 2044 19314 2096 19320
rect 2056 19009 2084 19314
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 2042 19000 2098 19009
rect 4214 19003 4522 19012
rect 2042 18935 2044 18944
rect 2096 18935 2098 18944
rect 2044 18906 2096 18912
rect 2056 18875 2084 18906
rect 1952 18760 2004 18766
rect 1952 18702 2004 18708
rect 1964 17882 1992 18702
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 2056 17785 2084 18226
rect 2042 17776 2098 17785
rect 2042 17711 2098 17720
rect 2044 16584 2096 16590
rect 1780 16546 1900 16574
rect 1492 16526 1544 16532
rect 1398 16416 1454 16425
rect 1398 16351 1454 16360
rect 1412 16114 1440 16351
rect 1504 16182 1532 16526
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 16250 1624 16390
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1492 16176 1544 16182
rect 1492 16118 1544 16124
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15858 1440 16050
rect 1412 15830 1532 15858
rect 1398 15736 1454 15745
rect 1504 15706 1532 15830
rect 1398 15671 1454 15680
rect 1492 15700 1544 15706
rect 1412 15502 1440 15671
rect 1492 15642 1544 15648
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1398 15328 1454 15337
rect 1398 15263 1454 15272
rect 1412 15042 1440 15263
rect 1412 15026 1532 15042
rect 1400 15020 1532 15026
rect 1452 15014 1532 15020
rect 1400 14962 1452 14968
rect 1398 14920 1454 14929
rect 1398 14855 1454 14864
rect 1412 14414 1440 14855
rect 1504 14618 1532 15014
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1596 14278 1624 14311
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1398 14104 1454 14113
rect 1398 14039 1454 14048
rect 1412 13938 1440 14039
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 12073 1440 12174
rect 1398 12064 1454 12073
rect 1454 12022 1532 12050
rect 1398 11999 1454 12008
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 1412 11150 1440 11591
rect 1504 11354 1532 12022
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1398 10840 1454 10849
rect 1398 10775 1454 10784
rect 1412 10674 1440 10775
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 9722 1440 10610
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10266 1624 10406
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1398 9616 1454 9625
rect 1398 9551 1400 9560
rect 1452 9551 1454 9560
rect 1400 9522 1452 9528
rect 1412 9330 1440 9522
rect 1412 9302 1532 9330
rect 1398 9208 1454 9217
rect 1504 9178 1532 9302
rect 1398 9143 1454 9152
rect 1492 9172 1544 9178
rect 1412 8974 1440 9143
rect 1492 9114 1544 9120
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8401 1440 8434
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 1412 8090 1440 8327
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1398 7984 1454 7993
rect 1398 7919 1454 7928
rect 1412 7886 1440 7919
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1780 7177 1808 7346
rect 1766 7168 1822 7177
rect 1766 7103 1822 7112
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1306 6352 1362 6361
rect 1306 6287 1362 6296
rect 1320 5234 1348 6287
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1504 5953 1532 6054
rect 1490 5944 1546 5953
rect 1490 5879 1546 5888
rect 1400 5636 1452 5642
rect 1400 5578 1452 5584
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1412 4146 1440 5578
rect 1780 5370 1808 6734
rect 1872 6662 1900 16546
rect 2044 16526 2096 16532
rect 2056 16153 2084 16526
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2042 16144 2098 16153
rect 2042 16079 2098 16088
rect 2240 15094 2268 16390
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2056 14521 2084 14962
rect 2042 14512 2098 14521
rect 2042 14447 2098 14456
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2056 13705 2084 13874
rect 2228 13728 2280 13734
rect 2042 13696 2098 13705
rect 2228 13670 2280 13676
rect 2042 13631 2098 13640
rect 2136 13320 2188 13326
rect 2134 13288 2136 13297
rect 2188 13288 2190 13297
rect 2134 13223 2190 13232
rect 2148 12442 2176 13223
rect 2240 12986 2268 13670
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2240 12481 2268 12718
rect 2226 12472 2282 12481
rect 2136 12436 2188 12442
rect 2226 12407 2228 12416
rect 2136 12378 2188 12384
rect 2280 12407 2282 12416
rect 2228 12378 2280 12384
rect 2240 12347 2268 12378
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11257 2268 11630
rect 2226 11248 2282 11257
rect 2226 11183 2282 11192
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 10441 2084 10610
rect 2042 10432 2098 10441
rect 2042 10367 2098 10376
rect 2228 10056 2280 10062
rect 2226 10024 2228 10033
rect 2280 10024 2282 10033
rect 2226 9959 2282 9968
rect 2332 8566 2360 18634
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 12918 2820 13262
rect 2780 12912 2832 12918
rect 2778 12880 2780 12889
rect 2832 12880 2834 12889
rect 2778 12815 2834 12824
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2332 8022 2360 8502
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 2780 6792 2832 6798
rect 2778 6760 2780 6769
rect 2832 6760 2834 6769
rect 2778 6695 2834 6704
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1872 5234 1900 6598
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1964 4826 1992 5578
rect 2148 5370 2176 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1964 3126 1992 4762
rect 2148 4214 2176 5306
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2792 4282 2820 5170
rect 3238 5128 3294 5137
rect 3238 5063 3294 5072
rect 3252 4622 3280 5063
rect 4632 5030 4660 22918
rect 13832 22642 13860 25434
rect 16592 23118 16620 26250
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 17788 20942 17816 24550
rect 19444 23730 19472 27270
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 37188 26308 37240 26314
rect 37188 26250 37240 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 37200 26042 37228 26250
rect 37188 26036 37240 26042
rect 37188 25978 37240 25984
rect 37188 25764 37240 25770
rect 37188 25706 37240 25712
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 37200 25498 37228 25706
rect 37188 25492 37240 25498
rect 37188 25434 37240 25440
rect 33140 25220 33192 25226
rect 33140 25162 33192 25168
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19800 24200 19852 24206
rect 19798 24168 19800 24177
rect 19852 24168 19854 24177
rect 19798 24103 19854 24112
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17880 20534 17908 22714
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13924 15434 13952 17206
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 14476 11762 14504 19722
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17880 17678 17908 19654
rect 17972 19514 18000 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21554 20024 24890
rect 33152 24818 33180 25162
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 37280 23520 37332 23526
rect 37280 23462 37332 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 37292 23322 37320 23462
rect 37280 23316 37332 23322
rect 37280 23258 37332 23264
rect 37292 23118 37320 23258
rect 37280 23112 37332 23118
rect 37280 23054 37332 23060
rect 31024 23044 31076 23050
rect 31024 22986 31076 22992
rect 31036 22642 31064 22986
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 37280 22432 37332 22438
rect 37280 22374 37332 22380
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 37292 22098 37320 22374
rect 37280 22092 37332 22098
rect 37280 22034 37332 22040
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 18972 20868 19024 20874
rect 18972 20810 19024 20816
rect 33140 20868 33192 20874
rect 33140 20810 33192 20816
rect 18984 20466 19012 20810
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 20466 19472 20742
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 33152 20602 33180 20810
rect 33140 20596 33192 20602
rect 33140 20538 33192 20544
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19168 20058 19196 20198
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18524 19718 18552 19790
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 15978 15148 16934
rect 17972 16590 18000 18090
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 15108 15972 15160 15978
rect 15108 15914 15160 15920
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15212 12238 15240 13126
rect 18432 12782 18460 19110
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13832 8906 13860 10202
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 15304 8634 15332 12106
rect 18524 10062 18552 19654
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 17066 18644 17478
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 19248 16584 19300 16590
rect 19444 16574 19472 20402
rect 19890 20360 19946 20369
rect 19890 20295 19892 20304
rect 19944 20295 19946 20304
rect 31024 20324 31076 20330
rect 19892 20266 19944 20272
rect 31024 20266 31076 20272
rect 21088 19984 21140 19990
rect 21088 19926 21140 19932
rect 20626 19816 20682 19825
rect 20626 19751 20628 19760
rect 20680 19751 20682 19760
rect 20628 19722 20680 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 21100 19378 21128 19926
rect 31036 19854 31064 20266
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 31760 20052 31812 20058
rect 31760 19994 31812 20000
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 27528 19508 27580 19514
rect 27528 19450 27580 19456
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20088 18086 20116 18702
rect 20364 18630 20392 19314
rect 21100 18970 21128 19314
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19248 16526 19300 16532
rect 19352 16546 19472 16574
rect 19260 16250 19288 16526
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19352 13394 19380 16546
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 13938 19472 14758
rect 19996 14414 20024 14826
rect 19984 14408 20036 14414
rect 20088 14385 20116 18022
rect 19984 14350 20036 14356
rect 20074 14376 20130 14385
rect 20074 14311 20130 14320
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 20364 14006 20392 18566
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20732 16794 20760 18090
rect 27540 17678 27568 19450
rect 31772 18970 31800 19994
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 31760 18964 31812 18970
rect 31760 18906 31812 18912
rect 37384 18630 37412 31334
rect 37476 19174 37504 33254
rect 37556 32768 37608 32774
rect 37556 32710 37608 32716
rect 37568 20369 37596 32710
rect 37648 30592 37700 30598
rect 37648 30534 37700 30540
rect 37554 20360 37610 20369
rect 37554 20295 37610 20304
rect 37660 19718 37688 30534
rect 37648 19712 37700 19718
rect 37648 19654 37700 19660
rect 37464 19168 37516 19174
rect 37464 19110 37516 19116
rect 37372 18624 37424 18630
rect 37372 18566 37424 18572
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 31036 17202 31064 17478
rect 31024 17196 31076 17202
rect 31024 17138 31076 17144
rect 37752 16998 37780 35634
rect 38016 35488 38068 35494
rect 38016 35430 38068 35436
rect 38028 35329 38056 35430
rect 38014 35320 38070 35329
rect 38014 35255 38070 35264
rect 38108 35080 38160 35086
rect 38108 35022 38160 35028
rect 38016 34944 38068 34950
rect 38016 34886 38068 34892
rect 38028 34649 38056 34886
rect 38014 34640 38070 34649
rect 38014 34575 38070 34584
rect 38014 33960 38070 33969
rect 38014 33895 38070 33904
rect 38028 33862 38056 33895
rect 38016 33856 38068 33862
rect 38016 33798 38068 33804
rect 38016 33312 38068 33318
rect 38014 33280 38016 33289
rect 38068 33280 38070 33289
rect 38014 33215 38070 33224
rect 38016 32768 38068 32774
rect 38016 32710 38068 32716
rect 38028 32609 38056 32710
rect 38014 32600 38070 32609
rect 38014 32535 38070 32544
rect 38016 32224 38068 32230
rect 38016 32166 38068 32172
rect 38028 31929 38056 32166
rect 38014 31920 38070 31929
rect 38014 31855 38070 31864
rect 37924 31340 37976 31346
rect 37924 31282 37976 31288
rect 37936 19825 37964 31282
rect 38014 31240 38070 31249
rect 38014 31175 38016 31184
rect 38068 31175 38070 31184
rect 38016 31146 38068 31152
rect 38016 30592 38068 30598
rect 38014 30560 38016 30569
rect 38068 30560 38070 30569
rect 38014 30495 38070 30504
rect 38016 30048 38068 30054
rect 38016 29990 38068 29996
rect 38028 29889 38056 29990
rect 38014 29880 38070 29889
rect 38014 29815 38070 29824
rect 38016 29504 38068 29510
rect 38016 29446 38068 29452
rect 38028 29209 38056 29446
rect 38014 29200 38070 29209
rect 38014 29135 38070 29144
rect 38014 28520 38070 28529
rect 38014 28455 38070 28464
rect 38028 28422 38056 28455
rect 38016 28416 38068 28422
rect 38016 28358 38068 28364
rect 38016 27872 38068 27878
rect 38014 27840 38016 27849
rect 38068 27840 38070 27849
rect 38014 27775 38070 27784
rect 38016 27328 38068 27334
rect 38016 27270 38068 27276
rect 38028 27169 38056 27270
rect 38014 27160 38070 27169
rect 38014 27095 38070 27104
rect 38016 26784 38068 26790
rect 38016 26726 38068 26732
rect 38028 26489 38056 26726
rect 38014 26480 38070 26489
rect 38014 26415 38070 26424
rect 38014 25800 38070 25809
rect 38014 25735 38016 25744
rect 38068 25735 38070 25744
rect 38016 25706 38068 25712
rect 38016 25152 38068 25158
rect 38014 25120 38016 25129
rect 38068 25120 38070 25129
rect 38014 25055 38070 25064
rect 38016 24608 38068 24614
rect 38016 24550 38068 24556
rect 38028 24449 38056 24550
rect 38014 24440 38070 24449
rect 38014 24375 38070 24384
rect 38016 24064 38068 24070
rect 38016 24006 38068 24012
rect 38028 23769 38056 24006
rect 38014 23760 38070 23769
rect 38014 23695 38070 23704
rect 38014 23080 38070 23089
rect 38014 23015 38070 23024
rect 38028 22982 38056 23015
rect 38016 22976 38068 22982
rect 38016 22918 38068 22924
rect 38016 22432 38068 22438
rect 38014 22400 38016 22409
rect 38068 22400 38070 22409
rect 38014 22335 38070 22344
rect 38016 21888 38068 21894
rect 38016 21830 38068 21836
rect 38028 21729 38056 21830
rect 38014 21720 38070 21729
rect 38014 21655 38070 21664
rect 38016 21344 38068 21350
rect 38016 21286 38068 21292
rect 38028 21049 38056 21286
rect 38014 21040 38070 21049
rect 38014 20975 38070 20984
rect 38014 20360 38070 20369
rect 38014 20295 38016 20304
rect 38068 20295 38070 20304
rect 38016 20266 38068 20272
rect 37922 19816 37978 19825
rect 37922 19751 37978 19760
rect 38016 19712 38068 19718
rect 38014 19680 38016 19689
rect 38068 19680 38070 19689
rect 38014 19615 38070 19624
rect 38016 19168 38068 19174
rect 38016 19110 38068 19116
rect 38028 19009 38056 19110
rect 38014 19000 38070 19009
rect 38014 18935 38070 18944
rect 38016 18624 38068 18630
rect 38016 18566 38068 18572
rect 38028 18329 38056 18566
rect 38014 18320 38070 18329
rect 38014 18255 38070 18264
rect 38014 17640 38070 17649
rect 38014 17575 38070 17584
rect 38028 17542 38056 17575
rect 38016 17536 38068 17542
rect 38016 17478 38068 17484
rect 38120 17066 38148 35022
rect 38212 17610 38240 36110
rect 38292 32428 38344 32434
rect 38292 32370 38344 32376
rect 38304 19242 38332 32370
rect 38292 19236 38344 19242
rect 38292 19178 38344 19184
rect 38200 17604 38252 17610
rect 38200 17546 38252 17552
rect 38108 17060 38160 17066
rect 38108 17002 38160 17008
rect 37740 16992 37792 16998
rect 38016 16992 38068 16998
rect 37740 16934 37792 16940
rect 38014 16960 38016 16969
rect 38068 16960 38070 16969
rect 34934 16892 35242 16901
rect 38014 16895 38070 16904
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 37188 16448 37240 16454
rect 37188 16390 37240 16396
rect 38016 16448 38068 16454
rect 38016 16390 38068 16396
rect 37200 16250 37228 16390
rect 38028 16289 38056 16390
rect 38014 16280 38070 16289
rect 37188 16244 37240 16250
rect 38014 16215 38070 16224
rect 37188 16186 37240 16192
rect 33140 15972 33192 15978
rect 33140 15914 33192 15920
rect 33152 15162 33180 15914
rect 38016 15904 38068 15910
rect 38016 15846 38068 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 38028 15609 38056 15846
rect 38014 15600 38070 15609
rect 38014 15535 38070 15544
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 37280 14952 37332 14958
rect 37280 14894 37332 14900
rect 38014 14920 38070 14929
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 37292 14618 37320 14894
rect 38014 14855 38016 14864
rect 38068 14855 38070 14864
rect 38016 14826 38068 14832
rect 37280 14612 37332 14618
rect 37280 14554 37332 14560
rect 37188 14272 37240 14278
rect 38016 14272 38068 14278
rect 37188 14214 37240 14220
rect 38014 14240 38016 14249
rect 38068 14240 38070 14249
rect 37200 14074 37228 14214
rect 38014 14175 38070 14184
rect 37188 14068 37240 14074
rect 37188 14010 37240 14016
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 37188 13864 37240 13870
rect 37188 13806 37240 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 37200 13530 37228 13806
rect 38016 13728 38068 13734
rect 38016 13670 38068 13676
rect 38028 13569 38056 13670
rect 38014 13560 38070 13569
rect 37188 13524 37240 13530
rect 38014 13495 38070 13504
rect 37188 13466 37240 13472
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 38016 13184 38068 13190
rect 38016 13126 38068 13132
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 38028 12889 38056 13126
rect 38014 12880 38070 12889
rect 38014 12815 38070 12824
rect 37004 12640 37056 12646
rect 37004 12582 37056 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 37016 12442 37044 12582
rect 37004 12436 37056 12442
rect 37004 12378 37056 12384
rect 38014 12200 38070 12209
rect 38014 12135 38070 12144
rect 38028 12102 38056 12135
rect 37188 12096 37240 12102
rect 37188 12038 37240 12044
rect 38016 12096 38068 12102
rect 38016 12038 38068 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 37200 11898 37228 12038
rect 37188 11892 37240 11898
rect 37188 11834 37240 11840
rect 38016 11552 38068 11558
rect 38014 11520 38016 11529
rect 38068 11520 38070 11529
rect 34934 11452 35242 11461
rect 38014 11455 38070 11464
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 38016 11280 38068 11286
rect 38016 11222 38068 11228
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 38028 10849 38056 11222
rect 38014 10840 38070 10849
rect 38014 10775 38070 10784
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19720 10062 19748 10474
rect 37280 10464 37332 10470
rect 37280 10406 37332 10412
rect 38016 10464 38068 10470
rect 38016 10406 38068 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 37292 9926 37320 10406
rect 38028 10169 38056 10406
rect 38014 10160 38070 10169
rect 38014 10095 38070 10104
rect 37280 9920 37332 9926
rect 37280 9862 37332 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 18432 8090 18460 9318
rect 19720 8974 19748 9522
rect 38014 9480 38070 9489
rect 38014 9415 38016 9424
rect 38068 9415 38070 9424
rect 38016 9386 38068 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19444 8430 19472 8774
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20640 8498 20668 8842
rect 37280 8832 37332 8838
rect 38016 8832 38068 8838
rect 37280 8774 37332 8780
rect 38014 8800 38016 8809
rect 38068 8800 38070 8809
rect 37292 8566 37320 8774
rect 38014 8735 38070 8744
rect 37280 8560 37332 8566
rect 37280 8502 37332 8508
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 37372 8492 37424 8498
rect 37372 8434 37424 8440
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18616 7546 18644 8366
rect 19444 7886 19472 8366
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 20640 7886 20668 8230
rect 21284 7886 21312 8230
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 19444 7410 19472 7822
rect 37384 7818 37412 8434
rect 38016 8356 38068 8362
rect 38016 8298 38068 8304
rect 38028 8129 38056 8298
rect 38014 8120 38070 8129
rect 38014 8055 38070 8064
rect 37372 7812 37424 7818
rect 37372 7754 37424 7760
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 20640 7410 20668 7686
rect 38028 7449 38056 7686
rect 38014 7440 38070 7449
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20628 7404 20680 7410
rect 38014 7375 38070 7384
rect 20628 7346 20680 7352
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19536 6798 19564 7142
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 20088 6322 20116 7346
rect 37832 7200 37884 7206
rect 37832 7142 37884 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 37844 6798 37872 7142
rect 37832 6792 37884 6798
rect 37832 6734 37884 6740
rect 38014 6760 38070 6769
rect 38014 6695 38070 6704
rect 38028 6662 38056 6695
rect 37832 6656 37884 6662
rect 37832 6598 37884 6604
rect 38016 6656 38068 6662
rect 38016 6598 38068 6604
rect 37844 6322 37872 6598
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 37832 6112 37884 6118
rect 38016 6112 38068 6118
rect 37832 6054 37884 6060
rect 38014 6080 38016 6089
rect 38068 6080 38070 6089
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 37844 5710 37872 6054
rect 38014 6015 38070 6024
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 38016 5568 38068 5574
rect 38016 5510 38068 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 38028 5409 38056 5510
rect 38014 5400 38070 5409
rect 38014 5335 38070 5344
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 38028 4729 38056 4966
rect 38014 4720 38070 4729
rect 38014 4655 38070 4664
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2136 4208 2188 4214
rect 2136 4150 2188 4156
rect 38106 4040 38162 4049
rect 38106 3975 38108 3984
rect 38160 3975 38162 3984
rect 38108 3946 38160 3952
rect 37372 3936 37424 3942
rect 37372 3878 37424 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2056 3194 2084 3470
rect 37384 3398 37412 3878
rect 38108 3528 38160 3534
rect 38108 3470 38160 3476
rect 37372 3392 37424 3398
rect 38120 3369 38148 3470
rect 37372 3334 37424 3340
rect 38106 3360 38162 3369
rect 19574 3292 19882 3301
rect 38106 3295 38162 3304
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 38014 36644 38070 36680
rect 38014 36624 38016 36644
rect 38016 36624 38068 36644
rect 38068 36624 38070 36644
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 1398 34856 1454 34912
rect 2226 34448 2282 34504
rect 1490 34040 1546 34096
rect 1306 33632 1362 33688
rect 1398 33224 1454 33280
rect 1582 32408 1638 32464
rect 1398 30776 1454 30832
rect 1490 30368 1546 30424
rect 1490 29144 1546 29200
rect 1306 28736 1362 28792
rect 1398 28328 1454 28384
rect 1766 31592 1822 31648
rect 2226 31184 2282 31240
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 2870 32852 2872 32872
rect 2872 32852 2924 32872
rect 2924 32852 2926 32872
rect 2870 32816 2926 32852
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 3054 32000 3110 32056
rect 2042 29960 2098 30016
rect 1582 27512 1638 27568
rect 1490 27104 1546 27160
rect 1398 26696 1454 26752
rect 1490 25472 1546 25528
rect 1398 25064 1454 25120
rect 1490 24248 1546 24304
rect 1398 23432 1454 23488
rect 1490 23024 1546 23080
rect 1398 22752 1454 22808
rect 1398 22208 1454 22264
rect 1398 21800 1454 21856
rect 1398 21392 1454 21448
rect 1490 21004 1546 21040
rect 1490 20984 1492 21004
rect 1492 20984 1544 21004
rect 1544 20984 1546 21004
rect 1398 19760 1454 19816
rect 1398 18536 1454 18592
rect 1490 18128 1546 18184
rect 1398 17312 1454 17368
rect 1398 16904 1454 16960
rect 2226 29588 2228 29608
rect 2228 29588 2280 29608
rect 2280 29588 2282 29608
rect 2226 29552 2282 29588
rect 2226 27920 2282 27976
rect 2042 25880 2098 25936
rect 2134 24656 2190 24712
rect 2594 27648 2650 27704
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 38014 35980 38016 36000
rect 38016 35980 38068 36000
rect 38068 35980 38070 36000
rect 38014 35944 38070 35980
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 2594 26288 2650 26344
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 2778 23840 2834 23896
rect 2226 20576 2282 20632
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 2870 20168 2926 20224
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 2778 19388 2780 19408
rect 2780 19388 2832 19408
rect 2832 19388 2834 19408
rect 2778 19352 2834 19388
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 2042 18964 2098 19000
rect 2042 18944 2044 18964
rect 2044 18944 2096 18964
rect 2096 18944 2098 18964
rect 2042 17720 2098 17776
rect 1398 16360 1454 16416
rect 1398 15680 1454 15736
rect 1398 15272 1454 15328
rect 1398 14864 1454 14920
rect 1582 14320 1638 14376
rect 1398 14048 1454 14104
rect 1398 12008 1454 12064
rect 1398 11600 1454 11656
rect 1398 10784 1454 10840
rect 1398 9580 1454 9616
rect 1398 9560 1400 9580
rect 1400 9560 1452 9580
rect 1452 9560 1454 9580
rect 1398 9152 1454 9208
rect 1398 8336 1454 8392
rect 1398 7928 1454 7984
rect 1766 7112 1822 7168
rect 1306 6296 1362 6352
rect 1490 5888 1546 5944
rect 2042 16088 2098 16144
rect 2042 14456 2098 14512
rect 2042 13640 2098 13696
rect 2134 13268 2136 13288
rect 2136 13268 2188 13288
rect 2188 13268 2190 13288
rect 2134 13232 2190 13268
rect 2226 12436 2282 12472
rect 2226 12416 2228 12436
rect 2228 12416 2280 12436
rect 2280 12416 2282 12436
rect 2226 11192 2282 11248
rect 2042 10376 2098 10432
rect 2226 10004 2228 10024
rect 2228 10004 2280 10024
rect 2280 10004 2282 10024
rect 2226 9968 2282 10004
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 2778 12860 2780 12880
rect 2780 12860 2832 12880
rect 2832 12860 2834 12880
rect 2778 12824 2834 12860
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2778 6740 2780 6760
rect 2780 6740 2832 6760
rect 2832 6740 2834 6760
rect 2778 6704 2834 6740
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 3238 5072 3294 5128
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19798 24148 19800 24168
rect 19800 24148 19852 24168
rect 19852 24148 19854 24168
rect 19798 24112 19854 24148
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19890 20324 19946 20360
rect 19890 20304 19892 20324
rect 19892 20304 19944 20324
rect 19944 20304 19946 20324
rect 20626 19780 20682 19816
rect 20626 19760 20628 19780
rect 20628 19760 20680 19780
rect 20680 19760 20682 19780
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20074 14320 20130 14376
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 37554 20304 37610 20360
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 38014 35264 38070 35320
rect 38014 34584 38070 34640
rect 38014 33904 38070 33960
rect 38014 33260 38016 33280
rect 38016 33260 38068 33280
rect 38068 33260 38070 33280
rect 38014 33224 38070 33260
rect 38014 32544 38070 32600
rect 38014 31864 38070 31920
rect 38014 31204 38070 31240
rect 38014 31184 38016 31204
rect 38016 31184 38068 31204
rect 38068 31184 38070 31204
rect 38014 30540 38016 30560
rect 38016 30540 38068 30560
rect 38068 30540 38070 30560
rect 38014 30504 38070 30540
rect 38014 29824 38070 29880
rect 38014 29144 38070 29200
rect 38014 28464 38070 28520
rect 38014 27820 38016 27840
rect 38016 27820 38068 27840
rect 38068 27820 38070 27840
rect 38014 27784 38070 27820
rect 38014 27104 38070 27160
rect 38014 26424 38070 26480
rect 38014 25764 38070 25800
rect 38014 25744 38016 25764
rect 38016 25744 38068 25764
rect 38068 25744 38070 25764
rect 38014 25100 38016 25120
rect 38016 25100 38068 25120
rect 38068 25100 38070 25120
rect 38014 25064 38070 25100
rect 38014 24384 38070 24440
rect 38014 23704 38070 23760
rect 38014 23024 38070 23080
rect 38014 22380 38016 22400
rect 38016 22380 38068 22400
rect 38068 22380 38070 22400
rect 38014 22344 38070 22380
rect 38014 21664 38070 21720
rect 38014 20984 38070 21040
rect 38014 20324 38070 20360
rect 38014 20304 38016 20324
rect 38016 20304 38068 20324
rect 38068 20304 38070 20324
rect 37922 19760 37978 19816
rect 38014 19660 38016 19680
rect 38016 19660 38068 19680
rect 38068 19660 38070 19680
rect 38014 19624 38070 19660
rect 38014 18944 38070 19000
rect 38014 18264 38070 18320
rect 38014 17584 38070 17640
rect 38014 16940 38016 16960
rect 38016 16940 38068 16960
rect 38068 16940 38070 16960
rect 38014 16904 38070 16940
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 38014 16224 38070 16280
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 38014 15544 38070 15600
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 38014 14884 38070 14920
rect 38014 14864 38016 14884
rect 38016 14864 38068 14884
rect 38068 14864 38070 14884
rect 38014 14220 38016 14240
rect 38016 14220 38068 14240
rect 38068 14220 38070 14240
rect 38014 14184 38070 14220
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 38014 13504 38070 13560
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 38014 12824 38070 12880
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 38014 12144 38070 12200
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 38014 11500 38016 11520
rect 38016 11500 38068 11520
rect 38068 11500 38070 11520
rect 38014 11464 38070 11500
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 38014 10784 38070 10840
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 38014 10104 38070 10160
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 38014 9444 38070 9480
rect 38014 9424 38016 9444
rect 38016 9424 38068 9444
rect 38068 9424 38070 9444
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 38014 8780 38016 8800
rect 38016 8780 38068 8800
rect 38068 8780 38070 8800
rect 38014 8744 38070 8780
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 38014 8064 38070 8120
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 38014 7384 38070 7440
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 38014 6704 38070 6760
rect 38014 6060 38016 6080
rect 38016 6060 38068 6080
rect 38068 6060 38070 6080
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 38014 6024 38070 6060
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 38014 5344 38070 5400
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 38014 4664 38070 4720
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 38106 4004 38162 4040
rect 38106 3984 38108 4004
rect 38108 3984 38160 4004
rect 38160 3984 38162 4004
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38106 3304 38162 3360
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 38009 36682 38075 36685
rect 39200 36682 40000 36712
rect 38009 36680 40000 36682
rect 38009 36624 38014 36680
rect 38070 36624 40000 36680
rect 38009 36622 40000 36624
rect 38009 36619 38075 36622
rect 39200 36592 40000 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 38009 36002 38075 36005
rect 39200 36002 40000 36032
rect 38009 36000 40000 36002
rect 38009 35944 38014 36000
rect 38070 35944 40000 36000
rect 38009 35942 40000 35944
rect 38009 35939 38075 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 39200 35912 40000 35942
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 38009 35322 38075 35325
rect 39200 35322 40000 35352
rect 38009 35320 40000 35322
rect 38009 35264 38014 35320
rect 38070 35264 40000 35320
rect 38009 35262 40000 35264
rect 38009 35259 38075 35262
rect 39200 35232 40000 35262
rect 0 34914 800 34944
rect 1393 34914 1459 34917
rect 0 34912 1459 34914
rect 0 34856 1398 34912
rect 1454 34856 1459 34912
rect 0 34854 1459 34856
rect 0 34824 800 34854
rect 1393 34851 1459 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38009 34642 38075 34645
rect 39200 34642 40000 34672
rect 38009 34640 40000 34642
rect 38009 34584 38014 34640
rect 38070 34584 40000 34640
rect 38009 34582 40000 34584
rect 38009 34579 38075 34582
rect 39200 34552 40000 34582
rect 0 34506 800 34536
rect 2221 34506 2287 34509
rect 0 34504 2287 34506
rect 0 34448 2226 34504
rect 2282 34448 2287 34504
rect 0 34446 2287 34448
rect 0 34416 800 34446
rect 2221 34443 2287 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 34098 800 34128
rect 1485 34098 1551 34101
rect 0 34096 1551 34098
rect 0 34040 1490 34096
rect 1546 34040 1551 34096
rect 0 34038 1551 34040
rect 0 34008 800 34038
rect 1485 34035 1551 34038
rect 38009 33962 38075 33965
rect 39200 33962 40000 33992
rect 38009 33960 40000 33962
rect 38009 33904 38014 33960
rect 38070 33904 40000 33960
rect 38009 33902 40000 33904
rect 38009 33899 38075 33902
rect 39200 33872 40000 33902
rect 19570 33760 19886 33761
rect 0 33690 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 1301 33690 1367 33693
rect 0 33688 1367 33690
rect 0 33632 1306 33688
rect 1362 33632 1367 33688
rect 0 33630 1367 33632
rect 0 33600 800 33630
rect 1301 33627 1367 33630
rect 0 33282 800 33312
rect 1393 33282 1459 33285
rect 0 33280 1459 33282
rect 0 33224 1398 33280
rect 1454 33224 1459 33280
rect 0 33222 1459 33224
rect 0 33192 800 33222
rect 1393 33219 1459 33222
rect 38009 33282 38075 33285
rect 39200 33282 40000 33312
rect 38009 33280 40000 33282
rect 38009 33224 38014 33280
rect 38070 33224 40000 33280
rect 38009 33222 40000 33224
rect 38009 33219 38075 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 39200 33192 40000 33222
rect 34930 33151 35246 33152
rect 0 32874 800 32904
rect 2865 32874 2931 32877
rect 0 32872 2931 32874
rect 0 32816 2870 32872
rect 2926 32816 2931 32872
rect 0 32814 2931 32816
rect 0 32784 800 32814
rect 2865 32811 2931 32814
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 38009 32602 38075 32605
rect 39200 32602 40000 32632
rect 38009 32600 40000 32602
rect 38009 32544 38014 32600
rect 38070 32544 40000 32600
rect 38009 32542 40000 32544
rect 38009 32539 38075 32542
rect 39200 32512 40000 32542
rect 0 32466 800 32496
rect 1577 32466 1643 32469
rect 0 32464 1643 32466
rect 0 32408 1582 32464
rect 1638 32408 1643 32464
rect 0 32406 1643 32408
rect 0 32376 800 32406
rect 1577 32403 1643 32406
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 3049 32058 3115 32061
rect 0 32056 3115 32058
rect 0 32000 3054 32056
rect 3110 32000 3115 32056
rect 0 31998 3115 32000
rect 0 31968 800 31998
rect 3049 31995 3115 31998
rect 38009 31922 38075 31925
rect 39200 31922 40000 31952
rect 38009 31920 40000 31922
rect 38009 31864 38014 31920
rect 38070 31864 40000 31920
rect 38009 31862 40000 31864
rect 38009 31859 38075 31862
rect 39200 31832 40000 31862
rect 0 31650 800 31680
rect 1761 31650 1827 31653
rect 0 31648 1827 31650
rect 0 31592 1766 31648
rect 1822 31592 1827 31648
rect 0 31590 1827 31592
rect 0 31560 800 31590
rect 1761 31587 1827 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 0 31242 800 31272
rect 2221 31242 2287 31245
rect 0 31240 2287 31242
rect 0 31184 2226 31240
rect 2282 31184 2287 31240
rect 0 31182 2287 31184
rect 0 31152 800 31182
rect 2221 31179 2287 31182
rect 38009 31242 38075 31245
rect 39200 31242 40000 31272
rect 38009 31240 40000 31242
rect 38009 31184 38014 31240
rect 38070 31184 40000 31240
rect 38009 31182 40000 31184
rect 38009 31179 38075 31182
rect 39200 31152 40000 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 0 30834 800 30864
rect 1393 30834 1459 30837
rect 0 30832 1459 30834
rect 0 30776 1398 30832
rect 1454 30776 1459 30832
rect 0 30774 1459 30776
rect 0 30744 800 30774
rect 1393 30771 1459 30774
rect 38009 30562 38075 30565
rect 39200 30562 40000 30592
rect 38009 30560 40000 30562
rect 38009 30504 38014 30560
rect 38070 30504 40000 30560
rect 38009 30502 40000 30504
rect 38009 30499 38075 30502
rect 19570 30496 19886 30497
rect 0 30426 800 30456
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 39200 30472 40000 30502
rect 19570 30431 19886 30432
rect 1485 30426 1551 30429
rect 0 30424 1551 30426
rect 0 30368 1490 30424
rect 1546 30368 1551 30424
rect 0 30366 1551 30368
rect 0 30336 800 30366
rect 1485 30363 1551 30366
rect 0 30018 800 30048
rect 2037 30018 2103 30021
rect 0 30016 2103 30018
rect 0 29960 2042 30016
rect 2098 29960 2103 30016
rect 0 29958 2103 29960
rect 0 29928 800 29958
rect 2037 29955 2103 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 38009 29882 38075 29885
rect 39200 29882 40000 29912
rect 38009 29880 40000 29882
rect 38009 29824 38014 29880
rect 38070 29824 40000 29880
rect 38009 29822 40000 29824
rect 38009 29819 38075 29822
rect 39200 29792 40000 29822
rect 0 29610 800 29640
rect 2221 29610 2287 29613
rect 0 29608 2287 29610
rect 0 29552 2226 29608
rect 2282 29552 2287 29608
rect 0 29550 2287 29552
rect 0 29520 800 29550
rect 2221 29547 2287 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 0 29202 800 29232
rect 1485 29202 1551 29205
rect 0 29200 1551 29202
rect 0 29144 1490 29200
rect 1546 29144 1551 29200
rect 0 29142 1551 29144
rect 0 29112 800 29142
rect 1485 29139 1551 29142
rect 38009 29202 38075 29205
rect 39200 29202 40000 29232
rect 38009 29200 40000 29202
rect 38009 29144 38014 29200
rect 38070 29144 40000 29200
rect 38009 29142 40000 29144
rect 38009 29139 38075 29142
rect 39200 29112 40000 29142
rect 4210 28864 4526 28865
rect 0 28794 800 28824
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 1301 28794 1367 28797
rect 0 28792 1367 28794
rect 0 28736 1306 28792
rect 1362 28736 1367 28792
rect 0 28734 1367 28736
rect 0 28704 800 28734
rect 1301 28731 1367 28734
rect 38009 28522 38075 28525
rect 39200 28522 40000 28552
rect 38009 28520 40000 28522
rect 38009 28464 38014 28520
rect 38070 28464 40000 28520
rect 38009 28462 40000 28464
rect 38009 28459 38075 28462
rect 39200 28432 40000 28462
rect 0 28386 800 28416
rect 1393 28386 1459 28389
rect 0 28384 1459 28386
rect 0 28328 1398 28384
rect 1454 28328 1459 28384
rect 0 28326 1459 28328
rect 0 28296 800 28326
rect 1393 28323 1459 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 0 27978 800 28008
rect 2221 27978 2287 27981
rect 0 27976 2287 27978
rect 0 27920 2226 27976
rect 2282 27920 2287 27976
rect 0 27918 2287 27920
rect 0 27888 800 27918
rect 2221 27915 2287 27918
rect 38009 27842 38075 27845
rect 39200 27842 40000 27872
rect 38009 27840 40000 27842
rect 38009 27784 38014 27840
rect 38070 27784 40000 27840
rect 38009 27782 40000 27784
rect 38009 27779 38075 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 39200 27752 40000 27782
rect 34930 27711 35246 27712
rect 2589 27708 2655 27709
rect 2589 27704 2636 27708
rect 2700 27706 2706 27708
rect 2589 27648 2594 27704
rect 2589 27644 2636 27648
rect 2700 27646 2746 27706
rect 2700 27644 2706 27646
rect 2589 27643 2655 27644
rect 0 27570 800 27600
rect 1577 27570 1643 27573
rect 0 27568 1643 27570
rect 0 27512 1582 27568
rect 1638 27512 1643 27568
rect 0 27510 1643 27512
rect 0 27480 800 27510
rect 1577 27507 1643 27510
rect 19570 27232 19886 27233
rect 0 27162 800 27192
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 1485 27162 1551 27165
rect 0 27160 1551 27162
rect 0 27104 1490 27160
rect 1546 27104 1551 27160
rect 0 27102 1551 27104
rect 0 27072 800 27102
rect 1485 27099 1551 27102
rect 38009 27162 38075 27165
rect 39200 27162 40000 27192
rect 38009 27160 40000 27162
rect 38009 27104 38014 27160
rect 38070 27104 40000 27160
rect 38009 27102 40000 27104
rect 38009 27099 38075 27102
rect 39200 27072 40000 27102
rect 0 26754 800 26784
rect 1393 26754 1459 26757
rect 0 26752 1459 26754
rect 0 26696 1398 26752
rect 1454 26696 1459 26752
rect 0 26694 1459 26696
rect 0 26664 800 26694
rect 1393 26691 1459 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 38009 26482 38075 26485
rect 39200 26482 40000 26512
rect 38009 26480 40000 26482
rect 38009 26424 38014 26480
rect 38070 26424 40000 26480
rect 38009 26422 40000 26424
rect 38009 26419 38075 26422
rect 39200 26392 40000 26422
rect 0 26346 800 26376
rect 2589 26346 2655 26349
rect 0 26344 2655 26346
rect 0 26288 2594 26344
rect 2650 26288 2655 26344
rect 0 26286 2655 26288
rect 0 26256 800 26286
rect 2589 26283 2655 26286
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 0 25938 800 25968
rect 2037 25938 2103 25941
rect 0 25936 2103 25938
rect 0 25880 2042 25936
rect 2098 25880 2103 25936
rect 0 25878 2103 25880
rect 0 25848 800 25878
rect 2037 25875 2103 25878
rect 38009 25802 38075 25805
rect 39200 25802 40000 25832
rect 38009 25800 40000 25802
rect 38009 25744 38014 25800
rect 38070 25744 40000 25800
rect 38009 25742 40000 25744
rect 38009 25739 38075 25742
rect 39200 25712 40000 25742
rect 4210 25600 4526 25601
rect 0 25530 800 25560
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 1485 25530 1551 25533
rect 0 25528 1551 25530
rect 0 25472 1490 25528
rect 1546 25472 1551 25528
rect 0 25470 1551 25472
rect 0 25440 800 25470
rect 1485 25467 1551 25470
rect 0 25122 800 25152
rect 1393 25122 1459 25125
rect 0 25120 1459 25122
rect 0 25064 1398 25120
rect 1454 25064 1459 25120
rect 0 25062 1459 25064
rect 0 25032 800 25062
rect 1393 25059 1459 25062
rect 38009 25122 38075 25125
rect 39200 25122 40000 25152
rect 38009 25120 40000 25122
rect 38009 25064 38014 25120
rect 38070 25064 40000 25120
rect 38009 25062 40000 25064
rect 38009 25059 38075 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 39200 25032 40000 25062
rect 19570 24991 19886 24992
rect 0 24714 800 24744
rect 2129 24714 2195 24717
rect 0 24712 2195 24714
rect 0 24656 2134 24712
rect 2190 24656 2195 24712
rect 0 24654 2195 24656
rect 0 24624 800 24654
rect 2129 24651 2195 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 38009 24442 38075 24445
rect 39200 24442 40000 24472
rect 38009 24440 40000 24442
rect 38009 24384 38014 24440
rect 38070 24384 40000 24440
rect 38009 24382 40000 24384
rect 38009 24379 38075 24382
rect 39200 24352 40000 24382
rect 0 24306 800 24336
rect 1485 24306 1551 24309
rect 0 24304 1551 24306
rect 0 24248 1490 24304
rect 1546 24248 1551 24304
rect 0 24246 1551 24248
rect 0 24216 800 24246
rect 1485 24243 1551 24246
rect 2630 24108 2636 24172
rect 2700 24170 2706 24172
rect 19793 24170 19859 24173
rect 2700 24168 19859 24170
rect 2700 24112 19798 24168
rect 19854 24112 19859 24168
rect 2700 24110 19859 24112
rect 2700 24108 2706 24110
rect 19793 24107 19859 24110
rect 19570 23968 19886 23969
rect 0 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 2773 23898 2839 23901
rect 0 23896 2839 23898
rect 0 23840 2778 23896
rect 2834 23840 2839 23896
rect 0 23838 2839 23840
rect 0 23808 800 23838
rect 2773 23835 2839 23838
rect 38009 23762 38075 23765
rect 39200 23762 40000 23792
rect 38009 23760 40000 23762
rect 38009 23704 38014 23760
rect 38070 23704 40000 23760
rect 38009 23702 40000 23704
rect 38009 23699 38075 23702
rect 39200 23672 40000 23702
rect 0 23490 800 23520
rect 1393 23490 1459 23493
rect 0 23488 1459 23490
rect 0 23432 1398 23488
rect 1454 23432 1459 23488
rect 0 23430 1459 23432
rect 0 23400 800 23430
rect 1393 23427 1459 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23082 800 23112
rect 1485 23082 1551 23085
rect 0 23080 1551 23082
rect 0 23024 1490 23080
rect 1546 23024 1551 23080
rect 0 23022 1551 23024
rect 0 22992 800 23022
rect 1485 23019 1551 23022
rect 38009 23082 38075 23085
rect 39200 23082 40000 23112
rect 38009 23080 40000 23082
rect 38009 23024 38014 23080
rect 38070 23024 40000 23080
rect 38009 23022 40000 23024
rect 38009 23019 38075 23022
rect 39200 22992 40000 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 1393 22810 1459 22813
rect 1350 22808 1459 22810
rect 1350 22752 1398 22808
rect 1454 22752 1459 22808
rect 1350 22747 1459 22752
rect 0 22674 800 22704
rect 1350 22674 1410 22747
rect 0 22614 1410 22674
rect 0 22584 800 22614
rect 38009 22402 38075 22405
rect 39200 22402 40000 22432
rect 38009 22400 40000 22402
rect 38009 22344 38014 22400
rect 38070 22344 40000 22400
rect 38009 22342 40000 22344
rect 38009 22339 38075 22342
rect 4210 22336 4526 22337
rect 0 22266 800 22296
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 39200 22312 40000 22342
rect 34930 22271 35246 22272
rect 1393 22266 1459 22269
rect 0 22264 1459 22266
rect 0 22208 1398 22264
rect 1454 22208 1459 22264
rect 0 22206 1459 22208
rect 0 22176 800 22206
rect 1393 22203 1459 22206
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 38009 21722 38075 21725
rect 39200 21722 40000 21752
rect 38009 21720 40000 21722
rect 38009 21664 38014 21720
rect 38070 21664 40000 21720
rect 38009 21662 40000 21664
rect 38009 21659 38075 21662
rect 39200 21632 40000 21662
rect 0 21450 800 21480
rect 1393 21450 1459 21453
rect 0 21448 1459 21450
rect 0 21392 1398 21448
rect 1454 21392 1459 21448
rect 0 21390 1459 21392
rect 0 21360 800 21390
rect 1393 21387 1459 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 0 21042 800 21072
rect 1485 21042 1551 21045
rect 0 21040 1551 21042
rect 0 20984 1490 21040
rect 1546 20984 1551 21040
rect 0 20982 1551 20984
rect 0 20952 800 20982
rect 1485 20979 1551 20982
rect 38009 21042 38075 21045
rect 39200 21042 40000 21072
rect 38009 21040 40000 21042
rect 38009 20984 38014 21040
rect 38070 20984 40000 21040
rect 38009 20982 40000 20984
rect 38009 20979 38075 20982
rect 39200 20952 40000 20982
rect 19570 20704 19886 20705
rect 0 20634 800 20664
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 2221 20634 2287 20637
rect 0 20632 2287 20634
rect 0 20576 2226 20632
rect 2282 20576 2287 20632
rect 0 20574 2287 20576
rect 0 20544 800 20574
rect 2221 20571 2287 20574
rect 19885 20362 19951 20365
rect 37549 20362 37615 20365
rect 19885 20360 37615 20362
rect 19885 20304 19890 20360
rect 19946 20304 37554 20360
rect 37610 20304 37615 20360
rect 19885 20302 37615 20304
rect 19885 20299 19951 20302
rect 37549 20299 37615 20302
rect 38009 20362 38075 20365
rect 39200 20362 40000 20392
rect 38009 20360 40000 20362
rect 38009 20304 38014 20360
rect 38070 20304 40000 20360
rect 38009 20302 40000 20304
rect 38009 20299 38075 20302
rect 39200 20272 40000 20302
rect 0 20226 800 20256
rect 2865 20226 2931 20229
rect 0 20224 2931 20226
rect 0 20168 2870 20224
rect 2926 20168 2931 20224
rect 0 20166 2931 20168
rect 0 20136 800 20166
rect 2865 20163 2931 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 0 19818 800 19848
rect 1393 19818 1459 19821
rect 0 19816 1459 19818
rect 0 19760 1398 19816
rect 1454 19760 1459 19816
rect 0 19758 1459 19760
rect 0 19728 800 19758
rect 1393 19755 1459 19758
rect 20621 19818 20687 19821
rect 37917 19818 37983 19821
rect 20621 19816 37983 19818
rect 20621 19760 20626 19816
rect 20682 19760 37922 19816
rect 37978 19760 37983 19816
rect 20621 19758 37983 19760
rect 20621 19755 20687 19758
rect 37917 19755 37983 19758
rect 38009 19682 38075 19685
rect 39200 19682 40000 19712
rect 38009 19680 40000 19682
rect 38009 19624 38014 19680
rect 38070 19624 40000 19680
rect 38009 19622 40000 19624
rect 38009 19619 38075 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 39200 19592 40000 19622
rect 19570 19551 19886 19552
rect 0 19410 800 19440
rect 2773 19410 2839 19413
rect 0 19408 2839 19410
rect 0 19352 2778 19408
rect 2834 19352 2839 19408
rect 0 19350 2839 19352
rect 0 19320 800 19350
rect 2773 19347 2839 19350
rect 4210 19072 4526 19073
rect 0 19002 800 19032
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 2037 19002 2103 19005
rect 0 19000 2103 19002
rect 0 18944 2042 19000
rect 2098 18944 2103 19000
rect 0 18942 2103 18944
rect 0 18912 800 18942
rect 2037 18939 2103 18942
rect 38009 19002 38075 19005
rect 39200 19002 40000 19032
rect 38009 19000 40000 19002
rect 38009 18944 38014 19000
rect 38070 18944 40000 19000
rect 38009 18942 40000 18944
rect 38009 18939 38075 18942
rect 39200 18912 40000 18942
rect 0 18594 800 18624
rect 1393 18594 1459 18597
rect 0 18592 1459 18594
rect 0 18536 1398 18592
rect 1454 18536 1459 18592
rect 0 18534 1459 18536
rect 0 18504 800 18534
rect 1393 18531 1459 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 38009 18322 38075 18325
rect 39200 18322 40000 18352
rect 38009 18320 40000 18322
rect 38009 18264 38014 18320
rect 38070 18264 40000 18320
rect 38009 18262 40000 18264
rect 38009 18259 38075 18262
rect 39200 18232 40000 18262
rect 0 18186 800 18216
rect 1485 18186 1551 18189
rect 0 18184 1551 18186
rect 0 18128 1490 18184
rect 1546 18128 1551 18184
rect 0 18126 1551 18128
rect 0 18096 800 18126
rect 1485 18123 1551 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 2037 17778 2103 17781
rect 0 17776 2103 17778
rect 0 17720 2042 17776
rect 2098 17720 2103 17776
rect 0 17718 2103 17720
rect 0 17688 800 17718
rect 2037 17715 2103 17718
rect 38009 17642 38075 17645
rect 39200 17642 40000 17672
rect 38009 17640 40000 17642
rect 38009 17584 38014 17640
rect 38070 17584 40000 17640
rect 38009 17582 40000 17584
rect 38009 17579 38075 17582
rect 39200 17552 40000 17582
rect 19570 17440 19886 17441
rect 0 17370 800 17400
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 1393 17370 1459 17373
rect 0 17368 1459 17370
rect 0 17312 1398 17368
rect 1454 17312 1459 17368
rect 0 17310 1459 17312
rect 0 17280 800 17310
rect 1393 17307 1459 17310
rect 0 16962 800 16992
rect 1393 16962 1459 16965
rect 0 16960 1459 16962
rect 0 16904 1398 16960
rect 1454 16904 1459 16960
rect 0 16902 1459 16904
rect 0 16872 800 16902
rect 1393 16899 1459 16902
rect 38009 16962 38075 16965
rect 39200 16962 40000 16992
rect 38009 16960 40000 16962
rect 38009 16904 38014 16960
rect 38070 16904 40000 16960
rect 38009 16902 40000 16904
rect 38009 16899 38075 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 39200 16872 40000 16902
rect 34930 16831 35246 16832
rect 0 16554 800 16584
rect 0 16494 1456 16554
rect 0 16464 800 16494
rect 1396 16421 1456 16494
rect 1393 16416 1459 16421
rect 1393 16360 1398 16416
rect 1454 16360 1459 16416
rect 1393 16355 1459 16360
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 38009 16282 38075 16285
rect 39200 16282 40000 16312
rect 38009 16280 40000 16282
rect 38009 16224 38014 16280
rect 38070 16224 40000 16280
rect 38009 16222 40000 16224
rect 38009 16219 38075 16222
rect 39200 16192 40000 16222
rect 0 16146 800 16176
rect 2037 16146 2103 16149
rect 0 16144 2103 16146
rect 0 16088 2042 16144
rect 2098 16088 2103 16144
rect 0 16086 2103 16088
rect 0 16056 800 16086
rect 2037 16083 2103 16086
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 38009 15602 38075 15605
rect 39200 15602 40000 15632
rect 38009 15600 40000 15602
rect 38009 15544 38014 15600
rect 38070 15544 40000 15600
rect 38009 15542 40000 15544
rect 38009 15539 38075 15542
rect 39200 15512 40000 15542
rect 0 15330 800 15360
rect 1393 15330 1459 15333
rect 0 15328 1459 15330
rect 0 15272 1398 15328
rect 1454 15272 1459 15328
rect 0 15270 1459 15272
rect 0 15240 800 15270
rect 1393 15267 1459 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 0 14922 800 14952
rect 1393 14922 1459 14925
rect 0 14920 1459 14922
rect 0 14864 1398 14920
rect 1454 14864 1459 14920
rect 0 14862 1459 14864
rect 0 14832 800 14862
rect 1393 14859 1459 14862
rect 38009 14922 38075 14925
rect 39200 14922 40000 14952
rect 38009 14920 40000 14922
rect 38009 14864 38014 14920
rect 38070 14864 40000 14920
rect 38009 14862 40000 14864
rect 38009 14859 38075 14862
rect 39200 14832 40000 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 0 14514 800 14544
rect 2037 14514 2103 14517
rect 0 14512 2103 14514
rect 0 14456 2042 14512
rect 2098 14456 2103 14512
rect 0 14454 2103 14456
rect 0 14424 800 14454
rect 2037 14451 2103 14454
rect 1577 14378 1643 14381
rect 20069 14378 20135 14381
rect 1577 14376 20135 14378
rect 1577 14320 1582 14376
rect 1638 14320 20074 14376
rect 20130 14320 20135 14376
rect 1577 14318 20135 14320
rect 1577 14315 1643 14318
rect 20069 14315 20135 14318
rect 38009 14242 38075 14245
rect 39200 14242 40000 14272
rect 38009 14240 40000 14242
rect 38009 14184 38014 14240
rect 38070 14184 40000 14240
rect 38009 14182 40000 14184
rect 38009 14179 38075 14182
rect 19570 14176 19886 14177
rect 0 14106 800 14136
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 39200 14152 40000 14182
rect 19570 14111 19886 14112
rect 1393 14106 1459 14109
rect 0 14104 1459 14106
rect 0 14048 1398 14104
rect 1454 14048 1459 14104
rect 0 14046 1459 14048
rect 0 14016 800 14046
rect 1393 14043 1459 14046
rect 0 13698 800 13728
rect 2037 13698 2103 13701
rect 0 13696 2103 13698
rect 0 13640 2042 13696
rect 2098 13640 2103 13696
rect 0 13638 2103 13640
rect 0 13608 800 13638
rect 2037 13635 2103 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 38009 13562 38075 13565
rect 39200 13562 40000 13592
rect 38009 13560 40000 13562
rect 38009 13504 38014 13560
rect 38070 13504 40000 13560
rect 38009 13502 40000 13504
rect 38009 13499 38075 13502
rect 39200 13472 40000 13502
rect 0 13290 800 13320
rect 2129 13290 2195 13293
rect 0 13288 2195 13290
rect 0 13232 2134 13288
rect 2190 13232 2195 13288
rect 0 13230 2195 13232
rect 0 13200 800 13230
rect 2129 13227 2195 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 0 12882 800 12912
rect 2773 12882 2839 12885
rect 0 12880 2839 12882
rect 0 12824 2778 12880
rect 2834 12824 2839 12880
rect 0 12822 2839 12824
rect 0 12792 800 12822
rect 2773 12819 2839 12822
rect 38009 12882 38075 12885
rect 39200 12882 40000 12912
rect 38009 12880 40000 12882
rect 38009 12824 38014 12880
rect 38070 12824 40000 12880
rect 38009 12822 40000 12824
rect 38009 12819 38075 12822
rect 39200 12792 40000 12822
rect 4210 12544 4526 12545
rect 0 12474 800 12504
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 2221 12474 2287 12477
rect 0 12472 2287 12474
rect 0 12416 2226 12472
rect 2282 12416 2287 12472
rect 0 12414 2287 12416
rect 0 12384 800 12414
rect 2221 12411 2287 12414
rect 38009 12202 38075 12205
rect 39200 12202 40000 12232
rect 38009 12200 40000 12202
rect 38009 12144 38014 12200
rect 38070 12144 40000 12200
rect 38009 12142 40000 12144
rect 38009 12139 38075 12142
rect 39200 12112 40000 12142
rect 0 12066 800 12096
rect 1393 12066 1459 12069
rect 0 12064 1459 12066
rect 0 12008 1398 12064
rect 1454 12008 1459 12064
rect 0 12006 1459 12008
rect 0 11976 800 12006
rect 1393 12003 1459 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 38009 11522 38075 11525
rect 39200 11522 40000 11552
rect 38009 11520 40000 11522
rect 38009 11464 38014 11520
rect 38070 11464 40000 11520
rect 38009 11462 40000 11464
rect 38009 11459 38075 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 39200 11432 40000 11462
rect 34930 11391 35246 11392
rect 0 11250 800 11280
rect 2221 11250 2287 11253
rect 0 11248 2287 11250
rect 0 11192 2226 11248
rect 2282 11192 2287 11248
rect 0 11190 2287 11192
rect 0 11160 800 11190
rect 2221 11187 2287 11190
rect 19570 10912 19886 10913
rect 0 10842 800 10872
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 1393 10842 1459 10845
rect 0 10840 1459 10842
rect 0 10784 1398 10840
rect 1454 10784 1459 10840
rect 0 10782 1459 10784
rect 0 10752 800 10782
rect 1393 10779 1459 10782
rect 38009 10842 38075 10845
rect 39200 10842 40000 10872
rect 38009 10840 40000 10842
rect 38009 10784 38014 10840
rect 38070 10784 40000 10840
rect 38009 10782 40000 10784
rect 38009 10779 38075 10782
rect 39200 10752 40000 10782
rect 0 10434 800 10464
rect 2037 10434 2103 10437
rect 0 10432 2103 10434
rect 0 10376 2042 10432
rect 2098 10376 2103 10432
rect 0 10374 2103 10376
rect 0 10344 800 10374
rect 2037 10371 2103 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 38009 10162 38075 10165
rect 39200 10162 40000 10192
rect 38009 10160 40000 10162
rect 38009 10104 38014 10160
rect 38070 10104 40000 10160
rect 38009 10102 40000 10104
rect 38009 10099 38075 10102
rect 39200 10072 40000 10102
rect 0 10026 800 10056
rect 2221 10026 2287 10029
rect 0 10024 2287 10026
rect 0 9968 2226 10024
rect 2282 9968 2287 10024
rect 0 9966 2287 9968
rect 0 9936 800 9966
rect 2221 9963 2287 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 38009 9482 38075 9485
rect 39200 9482 40000 9512
rect 38009 9480 40000 9482
rect 38009 9424 38014 9480
rect 38070 9424 40000 9480
rect 38009 9422 40000 9424
rect 38009 9419 38075 9422
rect 39200 9392 40000 9422
rect 4210 9280 4526 9281
rect 0 9210 800 9240
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 0 8712 800 8832
rect 38009 8802 38075 8805
rect 39200 8802 40000 8832
rect 38009 8800 40000 8802
rect 38009 8744 38014 8800
rect 38070 8744 40000 8800
rect 38009 8742 40000 8744
rect 38009 8739 38075 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 39200 8712 40000 8742
rect 19570 8671 19886 8672
rect 0 8394 800 8424
rect 1393 8394 1459 8397
rect 0 8392 1459 8394
rect 0 8336 1398 8392
rect 1454 8336 1459 8392
rect 0 8334 1459 8336
rect 0 8304 800 8334
rect 1393 8331 1459 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 38009 8122 38075 8125
rect 39200 8122 40000 8152
rect 38009 8120 40000 8122
rect 38009 8064 38014 8120
rect 38070 8064 40000 8120
rect 38009 8062 40000 8064
rect 38009 8059 38075 8062
rect 39200 8032 40000 8062
rect 0 7986 800 8016
rect 1393 7986 1459 7989
rect 0 7984 1459 7986
rect 0 7928 1398 7984
rect 1454 7928 1459 7984
rect 0 7926 1459 7928
rect 0 7896 800 7926
rect 1393 7923 1459 7926
rect 19570 7648 19886 7649
rect 0 7488 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 38009 7442 38075 7445
rect 39200 7442 40000 7472
rect 38009 7440 40000 7442
rect 38009 7384 38014 7440
rect 38070 7384 40000 7440
rect 38009 7382 40000 7384
rect 38009 7379 38075 7382
rect 39200 7352 40000 7382
rect 0 7170 800 7200
rect 1761 7170 1827 7173
rect 0 7168 1827 7170
rect 0 7112 1766 7168
rect 1822 7112 1827 7168
rect 0 7110 1827 7112
rect 0 7080 800 7110
rect 1761 7107 1827 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6762 800 6792
rect 2773 6762 2839 6765
rect 0 6760 2839 6762
rect 0 6704 2778 6760
rect 2834 6704 2839 6760
rect 0 6702 2839 6704
rect 0 6672 800 6702
rect 2773 6699 2839 6702
rect 38009 6762 38075 6765
rect 39200 6762 40000 6792
rect 38009 6760 40000 6762
rect 38009 6704 38014 6760
rect 38070 6704 40000 6760
rect 38009 6702 40000 6704
rect 38009 6699 38075 6702
rect 39200 6672 40000 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 0 6354 800 6384
rect 1301 6354 1367 6357
rect 0 6352 1367 6354
rect 0 6296 1306 6352
rect 1362 6296 1367 6352
rect 0 6294 1367 6296
rect 0 6264 800 6294
rect 1301 6291 1367 6294
rect 38009 6082 38075 6085
rect 39200 6082 40000 6112
rect 38009 6080 40000 6082
rect 38009 6024 38014 6080
rect 38070 6024 40000 6080
rect 38009 6022 40000 6024
rect 38009 6019 38075 6022
rect 4210 6016 4526 6017
rect 0 5946 800 5976
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 39200 5992 40000 6022
rect 34930 5951 35246 5952
rect 1485 5946 1551 5949
rect 0 5944 1551 5946
rect 0 5888 1490 5944
rect 1546 5888 1551 5944
rect 0 5886 1551 5888
rect 0 5856 800 5886
rect 1485 5883 1551 5886
rect 0 5448 800 5568
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 38009 5402 38075 5405
rect 39200 5402 40000 5432
rect 38009 5400 40000 5402
rect 38009 5344 38014 5400
rect 38070 5344 40000 5400
rect 38009 5342 40000 5344
rect 38009 5339 38075 5342
rect 39200 5312 40000 5342
rect 0 5130 800 5160
rect 3233 5130 3299 5133
rect 0 5128 3299 5130
rect 0 5072 3238 5128
rect 3294 5072 3299 5128
rect 0 5070 3299 5072
rect 0 5040 800 5070
rect 3233 5067 3299 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 38009 4722 38075 4725
rect 39200 4722 40000 4752
rect 38009 4720 40000 4722
rect 38009 4664 38014 4720
rect 38070 4664 40000 4720
rect 38009 4662 40000 4664
rect 38009 4659 38075 4662
rect 39200 4632 40000 4662
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 38101 4042 38167 4045
rect 39200 4042 40000 4072
rect 38101 4040 40000 4042
rect 38101 3984 38106 4040
rect 38162 3984 40000 4040
rect 38101 3982 40000 3984
rect 38101 3979 38167 3982
rect 39200 3952 40000 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 38101 3362 38167 3365
rect 39200 3362 40000 3392
rect 38101 3360 40000 3362
rect 38101 3304 38106 3360
rect 38162 3304 40000 3360
rect 38101 3302 40000 3304
rect 38101 3299 38167 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 39200 3272 40000 3302
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 2636 27704 2700 27708
rect 2636 27648 2650 27704
rect 2650 27648 2700 27704
rect 2636 27644 2700 27648
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 2636 24108 2700 24172
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 2635 27708 2701 27709
rect 2635 27644 2636 27708
rect 2700 27644 2701 27708
rect 2635 27643 2701 27644
rect 2638 24173 2698 27643
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 2635 24172 2701 24173
rect 2635 24108 2636 24172
rect 2700 24108 2701 24172
rect 2635 24107 2701 24108
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18768 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__B
timestamp 1649977179
transform 1 0 18032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__B
timestamp 1649977179
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1649977179
transform -1 0 20976 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__B
timestamp 1649977179
transform 1 0 20240 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1649977179
transform -1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__B
timestamp 1649977179
transform -1 0 19228 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1649977179
transform -1 0 21160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform -1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform -1 0 21252 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform 1 0 18400 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform -1 0 19596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform 1 0 18952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform -1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform -1 0 20516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform -1 0 20516 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform -1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform -1 0 20608 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform -1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform -1 0 20792 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform -1 0 20792 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform -1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform -1 0 20608 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform -1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform -1 0 19412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform -1 0 21160 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform -1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform -1 0 18032 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 21160 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 20792 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 20792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform -1 0 20976 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform -1 0 20976 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform -1 0 20792 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 20608 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform -1 0 20424 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 20424 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform -1 0 20608 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform -1 0 20700 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform -1 0 20700 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform -1 0 20792 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1649977179
transform -1 0 20884 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1649977179
transform -1 0 20792 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform -1 0 20700 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 2760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 2576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 3404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 2852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 2208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 2208 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 2760 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 2852 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 2208 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 2208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 2760 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 2208 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 2852 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 3956 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 2852 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 2208 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 2852 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 3680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 2668 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 2852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 2208 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 2852 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 2760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 2208 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 2760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 2852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 2208 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 2852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 3404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 2760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 2208 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 2208 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 2208 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 2760 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 3312 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 2760 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 2760 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 2760 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 2208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 2760 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 2760 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 2852 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 2760 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 2208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 3220 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 2760 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 2852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 2208 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 1564 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 2760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 2852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 2208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 2208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 2208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 2668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1649977179
transform -1 0 37444 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1649977179
transform -1 0 37444 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1649977179
transform -1 0 37444 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1649977179
transform -1 0 37444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1649977179
transform -1 0 37444 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1649977179
transform 1 0 37352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 1649977179
transform -1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1649977179
transform -1 0 37444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1649977179
transform -1 0 37444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1649977179
transform -1 0 37444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output85_A
timestamp 1649977179
transform 1 0 37260 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1649977179
transform 1 0 37260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1649977179
transform -1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1649977179
transform -1 0 37444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1649977179
transform 1 0 37260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1649977179
transform 1 0 37260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1649977179
transform -1 0 37444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output97_A
timestamp 1649977179
transform 1 0 37260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output98_A
timestamp 1649977179
transform -1 0 37444 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output100_A
timestamp 1649977179
transform 1 0 37260 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output101_A
timestamp 1649977179
transform -1 0 37444 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output102_A
timestamp 1649977179
transform 1 0 37260 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output103_A
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output105_A
timestamp 1649977179
transform -1 0 37444 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output107_A
timestamp 1649977179
transform -1 0 37444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output108_A
timestamp 1649977179
transform 1 0 37260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output109_A
timestamp 1649977179
transform 1 0 37260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output110_A
timestamp 1649977179
transform -1 0 37444 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1649977179
transform 1 0 37260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1649977179
transform -1 0 37444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1649977179
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1649977179
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1649977179
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1649977179
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_36
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1649977179
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_11
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1649977179
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_397
timestamp 1649977179
transform 1 0 37628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1649977179
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_19
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_31
timestamp 1649977179
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_43
timestamp 1649977179
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_396
timestamp 1649977179
transform 1 0 37536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1649977179
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_31
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_43
timestamp 1649977179
transform 1 0 5060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_55
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1649977179
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1649977179
transform 1 0 1656 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_395
timestamp 1649977179
transform 1 0 37444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1649977179
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_397
timestamp 1649977179
transform 1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1649977179
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_19
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_212
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1649977179
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_10
timestamp 1649977179
transform 1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_17
timestamp 1649977179
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1649977179
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_210
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_234
timestamp 1649977179
transform 1 0 22632 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1649977179
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_397
timestamp 1649977179
transform 1 0 37628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1649977179
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_17
timestamp 1649977179
transform 1 0 2668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1649977179
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1649977179
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1649977179
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_186
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_192
timestamp 1649977179
transform 1 0 18768 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_201
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_207
timestamp 1649977179
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1649977179
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1649977179
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp 1649977179
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_206
timestamp 1649977179
transform 1 0 20056 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1649977179
transform 1 0 20884 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_222
timestamp 1649977179
transform 1 0 21528 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_234
timestamp 1649977179
transform 1 0 22632 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_246
timestamp 1649977179
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_397
timestamp 1649977179
transform 1 0 37628 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1649977179
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_6
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_16
timestamp 1649977179
transform 1 0 2576 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_28
timestamp 1649977179
transform 1 0 3680 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_40
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_197
timestamp 1649977179
transform 1 0 19228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_206
timestamp 1649977179
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1649977179
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1649977179
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_12
timestamp 1649977179
transform 1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_18
timestamp 1649977179
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_199
timestamp 1649977179
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_207
timestamp 1649977179
transform 1 0 20148 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1649977179
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_216
timestamp 1649977179
transform 1 0 20976 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_228
timestamp 1649977179
transform 1 0 22080 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_240
timestamp 1649977179
transform 1 0 23184 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_395
timestamp 1649977179
transform 1 0 37444 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1649977179
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1649977179
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_12
timestamp 1649977179
transform 1 0 2208 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_24
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_36
timestamp 1649977179
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1649977179
transform 1 0 19596 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_211
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1649977179
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1649977179
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_205
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_211
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_223
timestamp 1649977179
transform 1 0 21620 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_235
timestamp 1649977179
transform 1 0 22724 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1649977179
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_6
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_19
timestamp 1649977179
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_31
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_395
timestamp 1649977179
transform 1 0 37444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1649977179
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp 1649977179
transform 1 0 1656 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_12
timestamp 1649977179
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1649977179
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1649977179
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_212
timestamp 1649977179
transform 1 0 20608 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_224
timestamp 1649977179
transform 1 0 21712 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_236
timestamp 1649977179
transform 1 0 22816 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_397
timestamp 1649977179
transform 1 0 37628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1649977179
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_19
timestamp 1649977179
transform 1 0 2852 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_31
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_395
timestamp 1649977179
transform 1 0 37444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1649977179
transform 1 0 38180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1649977179
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_12
timestamp 1649977179
transform 1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_18
timestamp 1649977179
transform 1 0 2760 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_206
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_212
timestamp 1649977179
transform 1 0 20608 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_224
timestamp 1649977179
transform 1 0 21712 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_236
timestamp 1649977179
transform 1 0 22816 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1649977179
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_395
timestamp 1649977179
transform 1 0 37444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1649977179
transform 1 0 38180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_19
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_31
timestamp 1649977179
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_201
timestamp 1649977179
transform 1 0 19596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_206
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_212
timestamp 1649977179
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1649977179
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_395
timestamp 1649977179
transform 1 0 37444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1649977179
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1649977179
transform 1 0 1656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_13
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_25
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_37
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1649977179
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1649977179
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp 1649977179
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1649977179
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_395
timestamp 1649977179
transform 1 0 37444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1649977179
transform 1 0 38180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_6
timestamp 1649977179
transform 1 0 1656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1649977179
transform 1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_208
timestamp 1649977179
transform 1 0 20240 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_214
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_226
timestamp 1649977179
transform 1 0 21896 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_238
timestamp 1649977179
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1649977179
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_395
timestamp 1649977179
transform 1 0 37444 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1649977179
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_6
timestamp 1649977179
transform 1 0 1656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_13
timestamp 1649977179
transform 1 0 2300 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_19
timestamp 1649977179
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_31
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1649977179
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 1649977179
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_395
timestamp 1649977179
transform 1 0 37444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1649977179
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1649977179
transform 1 0 1656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1649977179
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1649977179
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_12
timestamp 1649977179
transform 1 0 2208 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_24
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_36
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1649977179
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_199
timestamp 1649977179
transform 1 0 19412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_212
timestamp 1649977179
transform 1 0 20608 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_395
timestamp 1649977179
transform 1 0 37444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1649977179
transform 1 0 38180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_6
timestamp 1649977179
transform 1 0 1656 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_13
timestamp 1649977179
transform 1 0 2300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1649977179
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_215
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_227
timestamp 1649977179
transform 1 0 21988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_239
timestamp 1649977179
transform 1 0 23092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_395
timestamp 1649977179
transform 1 0 37444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1649977179
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 1649977179
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_18
timestamp 1649977179
transform 1 0 2760 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_30
timestamp 1649977179
transform 1 0 3864 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_42
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1649977179
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_204
timestamp 1649977179
transform 1 0 19872 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_212
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1649977179
transform 1 0 38180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_6
timestamp 1649977179
transform 1 0 1656 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_12
timestamp 1649977179
transform 1 0 2208 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1649977179
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_212
timestamp 1649977179
transform 1 0 20608 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_218
timestamp 1649977179
transform 1 0 21160 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_230
timestamp 1649977179
transform 1 0 22264 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_242
timestamp 1649977179
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1649977179
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_395
timestamp 1649977179
transform 1 0 37444 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1649977179
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_6
timestamp 1649977179
transform 1 0 1656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1649977179
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_19
timestamp 1649977179
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1649977179
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1649977179
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_10
timestamp 1649977179
transform 1 0 2024 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_16
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_205
timestamp 1649977179
transform 1 0 19964 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_211
timestamp 1649977179
transform 1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_217
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_229
timestamp 1649977179
transform 1 0 22172 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1649977179
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1649977179
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_395
timestamp 1649977179
transform 1 0 37444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1649977179
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_6
timestamp 1649977179
transform 1 0 1656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_25
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_37
timestamp 1649977179
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1649977179
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1649977179
transform 1 0 18032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_190
timestamp 1649977179
transform 1 0 18584 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_213
timestamp 1649977179
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_395
timestamp 1649977179
transform 1 0 37444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1649977179
transform 1 0 38180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_14
timestamp 1649977179
transform 1 0 2392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1649977179
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_205
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_219
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_231
timestamp 1649977179
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1649977179
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_397
timestamp 1649977179
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1649977179
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_12
timestamp 1649977179
transform 1 0 2208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_19
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_25
timestamp 1649977179
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_37
timestamp 1649977179
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1649977179
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_212
timestamp 1649977179
transform 1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1649977179
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_395
timestamp 1649977179
transform 1 0 37444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1649977179
transform 1 0 38180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_6
timestamp 1649977179
transform 1 0 1656 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1649977179
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1649977179
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1649977179
transform 1 0 19596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1649977179
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_214
timestamp 1649977179
transform 1 0 20792 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_226
timestamp 1649977179
transform 1 0 21896 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_238
timestamp 1649977179
transform 1 0 23000 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1649977179
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_6
timestamp 1649977179
transform 1 0 1656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_12
timestamp 1649977179
transform 1 0 2208 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_18
timestamp 1649977179
transform 1 0 2760 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_30
timestamp 1649977179
transform 1 0 3864 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_42
timestamp 1649977179
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1649977179
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1649977179
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1649977179
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1649977179
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1649977179
transform 1 0 38180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_6
timestamp 1649977179
transform 1 0 1656 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_12
timestamp 1649977179
transform 1 0 2208 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_395
timestamp 1649977179
transform 1 0 37444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1649977179
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_6
timestamp 1649977179
transform 1 0 1656 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_12
timestamp 1649977179
transform 1 0 2208 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_24
timestamp 1649977179
transform 1 0 3312 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_36
timestamp 1649977179
transform 1 0 4416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1649977179
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_210
timestamp 1649977179
transform 1 0 20424 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1649977179
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1649977179
transform 1 0 38180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_6
timestamp 1649977179
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_12
timestamp 1649977179
transform 1 0 2208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_18
timestamp 1649977179
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1649977179
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_37
timestamp 1649977179
transform 1 0 4508 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_49
timestamp 1649977179
transform 1 0 5612 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_61
timestamp 1649977179
transform 1 0 6716 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_73
timestamp 1649977179
transform 1 0 7820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_81
timestamp 1649977179
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_205
timestamp 1649977179
transform 1 0 19964 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1649977179
transform 1 0 20424 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_216
timestamp 1649977179
transform 1 0 20976 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_228
timestamp 1649977179
transform 1 0 22080 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_240
timestamp 1649977179
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_395
timestamp 1649977179
transform 1 0 37444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1649977179
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_6
timestamp 1649977179
transform 1 0 1656 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_18
timestamp 1649977179
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_30
timestamp 1649977179
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_42
timestamp 1649977179
transform 1 0 4968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1649977179
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_208
timestamp 1649977179
transform 1 0 20240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_214
timestamp 1649977179
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1649977179
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_12
timestamp 1649977179
transform 1 0 2208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_19
timestamp 1649977179
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_206
timestamp 1649977179
transform 1 0 20056 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_212
timestamp 1649977179
transform 1 0 20608 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_224
timestamp 1649977179
transform 1 0 21712 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_236
timestamp 1649977179
transform 1 0 22816 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1649977179
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_397
timestamp 1649977179
transform 1 0 37628 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1649977179
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_6
timestamp 1649977179
transform 1 0 1656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_13
timestamp 1649977179
transform 1 0 2300 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1649977179
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1649977179
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1649977179
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_395
timestamp 1649977179
transform 1 0 37444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1649977179
transform 1 0 38180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_6
timestamp 1649977179
transform 1 0 1656 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_12
timestamp 1649977179
transform 1 0 2208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_18
timestamp 1649977179
transform 1 0 2760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1649977179
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_204
timestamp 1649977179
transform 1 0 19872 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_210
timestamp 1649977179
transform 1 0 20424 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_222
timestamp 1649977179
transform 1 0 21528 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_234
timestamp 1649977179
transform 1 0 22632 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_246
timestamp 1649977179
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_395
timestamp 1649977179
transform 1 0 37444 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 1649977179
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_6
timestamp 1649977179
transform 1 0 1656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_12
timestamp 1649977179
transform 1 0 2208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_18
timestamp 1649977179
transform 1 0 2760 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_24
timestamp 1649977179
transform 1 0 3312 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_36
timestamp 1649977179
transform 1 0 4416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_48
timestamp 1649977179
transform 1 0 5520 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_204
timestamp 1649977179
transform 1 0 19872 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_210
timestamp 1649977179
transform 1 0 20424 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1649977179
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_395
timestamp 1649977179
transform 1 0 37444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1649977179
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_6
timestamp 1649977179
transform 1 0 1656 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_13
timestamp 1649977179
transform 1 0 2300 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1649977179
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1649977179
transform 1 0 20056 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_212
timestamp 1649977179
transform 1 0 20608 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_224
timestamp 1649977179
transform 1 0 21712 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_236
timestamp 1649977179
transform 1 0 22816 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1649977179
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_12
timestamp 1649977179
transform 1 0 2208 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_18
timestamp 1649977179
transform 1 0 2760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_30
timestamp 1649977179
transform 1 0 3864 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_42
timestamp 1649977179
transform 1 0 4968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1649977179
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_201
timestamp 1649977179
transform 1 0 19596 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_207
timestamp 1649977179
transform 1 0 20148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_213
timestamp 1649977179
transform 1 0 20700 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1649977179
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1649977179
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1649977179
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_12
timestamp 1649977179
transform 1 0 2208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_18
timestamp 1649977179
transform 1 0 2760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1649977179
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_395
timestamp 1649977179
transform 1 0 37444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1649977179
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_6
timestamp 1649977179
transform 1 0 1656 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_13
timestamp 1649977179
transform 1 0 2300 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_19
timestamp 1649977179
transform 1 0 2852 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_31
timestamp 1649977179
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1649977179
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_201
timestamp 1649977179
transform 1 0 19596 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_207
timestamp 1649977179
transform 1 0 20148 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1649977179
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1649977179
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_395
timestamp 1649977179
transform 1 0 37444 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1649977179
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_6
timestamp 1649977179
transform 1 0 1656 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_12
timestamp 1649977179
transform 1 0 2208 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1649977179
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1649977179
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_214
timestamp 1649977179
transform 1 0 20792 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_226
timestamp 1649977179
transform 1 0 21896 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_238
timestamp 1649977179
transform 1 0 23000 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1649977179
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_395
timestamp 1649977179
transform 1 0 37444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1649977179
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_6
timestamp 1649977179
transform 1 0 1656 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_12
timestamp 1649977179
transform 1 0 2208 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_18
timestamp 1649977179
transform 1 0 2760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_30
timestamp 1649977179
transform 1 0 3864 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_42
timestamp 1649977179
transform 1 0 4968 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1649977179
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_209
timestamp 1649977179
transform 1 0 20332 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_215
timestamp 1649977179
transform 1 0 20884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1649977179
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_6
timestamp 1649977179
transform 1 0 1656 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_13
timestamp 1649977179
transform 1 0 2300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_31
timestamp 1649977179
transform 1 0 3956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_43
timestamp 1649977179
transform 1 0 5060 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_55
timestamp 1649977179
transform 1 0 6164 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_67
timestamp 1649977179
transform 1 0 7268 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_79
timestamp 1649977179
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1649977179
transform 1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_214
timestamp 1649977179
transform 1 0 20792 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_226
timestamp 1649977179
transform 1 0 21896 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_238
timestamp 1649977179
transform 1 0 23000 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1649977179
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_397
timestamp 1649977179
transform 1 0 37628 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1649977179
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_6
timestamp 1649977179
transform 1 0 1656 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_13
timestamp 1649977179
transform 1 0 2300 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_19
timestamp 1649977179
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1649977179
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1649977179
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_395
timestamp 1649977179
transform 1 0 37444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1649977179
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_12
timestamp 1649977179
transform 1 0 2208 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_18
timestamp 1649977179
transform 1 0 2760 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1649977179
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_203
timestamp 1649977179
transform 1 0 19780 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_207
timestamp 1649977179
transform 1 0 20148 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_213
timestamp 1649977179
transform 1 0 20700 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_225
timestamp 1649977179
transform 1 0 21804 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_237
timestamp 1649977179
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1649977179
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_395
timestamp 1649977179
transform 1 0 37444 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1649977179
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_6
timestamp 1649977179
transform 1 0 1656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_13
timestamp 1649977179
transform 1 0 2300 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_19
timestamp 1649977179
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_31
timestamp 1649977179
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_43
timestamp 1649977179
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_395
timestamp 1649977179
transform 1 0 37444 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1649977179
transform 1 0 38180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_6
timestamp 1649977179
transform 1 0 1656 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_12
timestamp 1649977179
transform 1 0 2208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_18
timestamp 1649977179
transform 1 0 2760 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1649977179
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_6
timestamp 1649977179
transform 1 0 1656 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_22
timestamp 1649977179
transform 1 0 3128 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_28
timestamp 1649977179
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_40
timestamp 1649977179
transform 1 0 4784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1649977179
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_395
timestamp 1649977179
transform 1 0 37444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1649977179
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_13
timestamp 1649977179
transform 1 0 2300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1649977179
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_395
timestamp 1649977179
transform 1 0 37444 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1649977179
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_6
timestamp 1649977179
transform 1 0 1656 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_14
timestamp 1649977179
transform 1 0 2392 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_17
timestamp 1649977179
transform 1 0 2668 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_23
timestamp 1649977179
transform 1 0 3220 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_35
timestamp 1649977179
transform 1 0 4324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 1649977179
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_395
timestamp 1649977179
transform 1 0 37444 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1649977179
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_6
timestamp 1649977179
transform 1 0 1656 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_12
timestamp 1649977179
transform 1 0 2208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1649977179
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1649977179
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_395
timestamp 1649977179
transform 1 0 37444 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1649977179
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_6
timestamp 1649977179
transform 1 0 1656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_13
timestamp 1649977179
transform 1 0 2300 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_19
timestamp 1649977179
transform 1 0 2852 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_31
timestamp 1649977179
transform 1 0 3956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_43
timestamp 1649977179
transform 1 0 5060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_6
timestamp 1649977179
transform 1 0 1656 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_12
timestamp 1649977179
transform 1 0 2208 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1649977179
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_395
timestamp 1649977179
transform 1 0 37444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1649977179
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_6
timestamp 1649977179
transform 1 0 1656 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_12
timestamp 1649977179
transform 1 0 2208 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_24
timestamp 1649977179
transform 1 0 3312 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_36
timestamp 1649977179
transform 1 0 4416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_48
timestamp 1649977179
transform 1 0 5520 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_395
timestamp 1649977179
transform 1 0 37444 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1649977179
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_5
timestamp 1649977179
transform 1 0 1564 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_17
timestamp 1649977179
transform 1 0 2668 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_25
timestamp 1649977179
transform 1 0 3404 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_395
timestamp 1649977179
transform 1 0 37444 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1649977179
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_395
timestamp 1649977179
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1649977179
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_57
timestamp 1649977179
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_69
timestamp 1649977179
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1649977179
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1649977179
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1649977179
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1649977179
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_169
timestamp 1649977179
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_181
timestamp 1649977179
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1649977179
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_225
timestamp 1649977179
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1649977179
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1649977179
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_281
timestamp 1649977179
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_293
timestamp 1649977179
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1649977179
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_337
timestamp 1649977179
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_349
timestamp 1649977179
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1649977179
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_393
timestamp 1649977179
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1649977179
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _13_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _14_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _15_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _16_
timestamp 1649977179
transform 1 0 1840 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _17_
timestamp 1649977179
transform 1 0 1656 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _18_
timestamp 1649977179
transform 1 0 1656 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _19_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _20_
timestamp 1649977179
transform -1 0 2208 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _21_
timestamp 1649977179
transform 1 0 2208 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _22_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _23_
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _24_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2024 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _25_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19136 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _26_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _27_
timestamp 1649977179
transform 1 0 19596 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1649977179
transform -1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _29_
timestamp 1649977179
transform 1 0 20424 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1649977179
transform -1 0 21528 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _31_
timestamp 1649977179
transform 1 0 19596 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1649977179
transform -1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _33_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _34_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _36_
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _37_
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _38_
timestamp 1649977179
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _39_
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _40_
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _41_
timestamp 1649977179
transform 1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _42_
timestamp 1649977179
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _43_
timestamp 1649977179
transform 1 0 19504 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _44_
timestamp 1649977179
transform 1 0 19596 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_ pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _46_
timestamp 1649977179
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform -1 0 19964 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform -1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform -1 0 20056 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform -1 0 20056 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform -1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform -1 0 20240 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform -1 0 20240 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform -1 0 20240 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 20056 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 19688 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 20608 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform -1 0 21344 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 19228 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform -1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform -1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform -1 0 20240 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 20240 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 20424 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 20424 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 20240 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 20056 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 19872 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 19872 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 20056 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform -1 0 20148 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform -1 0 20148 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform -1 0 20240 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform -1 0 20332 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform -1 0 20240 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform -1 0 20148 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1649977179
transform -1 0 3312 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 1656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 2576 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 2668 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 1656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 2024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 1656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 1656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 2024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 2852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform 1 0 2668 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 1656 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 2024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 2300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 2852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform -1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 2300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform -1 0 1656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform -1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform -1 0 1656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform -1 0 2300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform -1 0 1656 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform -1 0 1656 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform -1 0 2300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform -1 0 1656 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform -1 0 1656 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 2944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 2300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 2300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1649977179
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1649977179
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform 1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 37812 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 37812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 37812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 37812 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 37812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 37812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 37812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 37812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 37812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output79
timestamp 1649977179
transform -1 0 38180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 37812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 37812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 37812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 37812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 37812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 37812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 37812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 37812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 37812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 37812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 37812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 37812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 37812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 37812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 37812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 37812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 37812 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 37812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 37812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 37812 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 37812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 37812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform 1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 37812 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 37812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform 1 0 37812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 37812 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 37812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 37812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 37812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  wb_interface_120 pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37904 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal3 s 39200 30472 40000 30592 0 FreeSans 480 0 0 0 addr0[0]
port 0 nsew signal tristate
flabel metal3 s 39200 31152 40000 31272 0 FreeSans 480 0 0 0 addr0[1]
port 1 nsew signal tristate
flabel metal3 s 39200 31832 40000 31952 0 FreeSans 480 0 0 0 addr0[2]
port 2 nsew signal tristate
flabel metal3 s 39200 32512 40000 32632 0 FreeSans 480 0 0 0 addr0[3]
port 3 nsew signal tristate
flabel metal3 s 39200 33192 40000 33312 0 FreeSans 480 0 0 0 addr0[4]
port 4 nsew signal tristate
flabel metal3 s 39200 33872 40000 33992 0 FreeSans 480 0 0 0 addr0[5]
port 5 nsew signal tristate
flabel metal3 s 39200 34552 40000 34672 0 FreeSans 480 0 0 0 addr0[6]
port 6 nsew signal tristate
flabel metal3 s 39200 35232 40000 35352 0 FreeSans 480 0 0 0 addr0[7]
port 7 nsew signal tristate
flabel metal3 s 39200 35912 40000 36032 0 FreeSans 480 0 0 0 addr0[8]
port 8 nsew signal tristate
flabel metal3 s 39200 3952 40000 4072 0 FreeSans 480 0 0 0 clk0
port 9 nsew signal tristate
flabel metal3 s 39200 4632 40000 4752 0 FreeSans 480 0 0 0 csb0
port 10 nsew signal tristate
flabel metal3 s 39200 8712 40000 8832 0 FreeSans 480 0 0 0 din0[0]
port 11 nsew signal tristate
flabel metal3 s 39200 15512 40000 15632 0 FreeSans 480 0 0 0 din0[10]
port 12 nsew signal tristate
flabel metal3 s 39200 16192 40000 16312 0 FreeSans 480 0 0 0 din0[11]
port 13 nsew signal tristate
flabel metal3 s 39200 16872 40000 16992 0 FreeSans 480 0 0 0 din0[12]
port 14 nsew signal tristate
flabel metal3 s 39200 17552 40000 17672 0 FreeSans 480 0 0 0 din0[13]
port 15 nsew signal tristate
flabel metal3 s 39200 18232 40000 18352 0 FreeSans 480 0 0 0 din0[14]
port 16 nsew signal tristate
flabel metal3 s 39200 18912 40000 19032 0 FreeSans 480 0 0 0 din0[15]
port 17 nsew signal tristate
flabel metal3 s 39200 19592 40000 19712 0 FreeSans 480 0 0 0 din0[16]
port 18 nsew signal tristate
flabel metal3 s 39200 20272 40000 20392 0 FreeSans 480 0 0 0 din0[17]
port 19 nsew signal tristate
flabel metal3 s 39200 20952 40000 21072 0 FreeSans 480 0 0 0 din0[18]
port 20 nsew signal tristate
flabel metal3 s 39200 21632 40000 21752 0 FreeSans 480 0 0 0 din0[19]
port 21 nsew signal tristate
flabel metal3 s 39200 9392 40000 9512 0 FreeSans 480 0 0 0 din0[1]
port 22 nsew signal tristate
flabel metal3 s 39200 22312 40000 22432 0 FreeSans 480 0 0 0 din0[20]
port 23 nsew signal tristate
flabel metal3 s 39200 22992 40000 23112 0 FreeSans 480 0 0 0 din0[21]
port 24 nsew signal tristate
flabel metal3 s 39200 23672 40000 23792 0 FreeSans 480 0 0 0 din0[22]
port 25 nsew signal tristate
flabel metal3 s 39200 24352 40000 24472 0 FreeSans 480 0 0 0 din0[23]
port 26 nsew signal tristate
flabel metal3 s 39200 25032 40000 25152 0 FreeSans 480 0 0 0 din0[24]
port 27 nsew signal tristate
flabel metal3 s 39200 25712 40000 25832 0 FreeSans 480 0 0 0 din0[25]
port 28 nsew signal tristate
flabel metal3 s 39200 26392 40000 26512 0 FreeSans 480 0 0 0 din0[26]
port 29 nsew signal tristate
flabel metal3 s 39200 27072 40000 27192 0 FreeSans 480 0 0 0 din0[27]
port 30 nsew signal tristate
flabel metal3 s 39200 27752 40000 27872 0 FreeSans 480 0 0 0 din0[28]
port 31 nsew signal tristate
flabel metal3 s 39200 28432 40000 28552 0 FreeSans 480 0 0 0 din0[29]
port 32 nsew signal tristate
flabel metal3 s 39200 10072 40000 10192 0 FreeSans 480 0 0 0 din0[2]
port 33 nsew signal tristate
flabel metal3 s 39200 29112 40000 29232 0 FreeSans 480 0 0 0 din0[30]
port 34 nsew signal tristate
flabel metal3 s 39200 29792 40000 29912 0 FreeSans 480 0 0 0 din0[31]
port 35 nsew signal tristate
flabel metal3 s 39200 10752 40000 10872 0 FreeSans 480 0 0 0 din0[3]
port 36 nsew signal tristate
flabel metal3 s 39200 11432 40000 11552 0 FreeSans 480 0 0 0 din0[4]
port 37 nsew signal tristate
flabel metal3 s 39200 12112 40000 12232 0 FreeSans 480 0 0 0 din0[5]
port 38 nsew signal tristate
flabel metal3 s 39200 12792 40000 12912 0 FreeSans 480 0 0 0 din0[6]
port 39 nsew signal tristate
flabel metal3 s 39200 13472 40000 13592 0 FreeSans 480 0 0 0 din0[7]
port 40 nsew signal tristate
flabel metal3 s 39200 14152 40000 14272 0 FreeSans 480 0 0 0 din0[8]
port 41 nsew signal tristate
flabel metal3 s 39200 14832 40000 14952 0 FreeSans 480 0 0 0 din0[9]
port 42 nsew signal tristate
flabel metal3 s 39200 3272 40000 3392 0 FreeSans 480 0 0 0 imem_rd_cs1
port 43 nsew signal tristate
flabel metal3 s 39200 36592 40000 36712 0 FreeSans 480 0 0 0 processor_reset
port 44 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 45 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 45 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 46 nsew ground bidirectional
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 wb_clk_i
port 47 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 wb_rst_i
port 48 nsew signal input
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 wbs_ack_o
port 49 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 wbs_adr_i[0]
port 50 nsew signal input
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 wbs_adr_i[10]
port 51 nsew signal input
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 wbs_adr_i[11]
port 52 nsew signal input
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 wbs_adr_i[12]
port 53 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 wbs_adr_i[13]
port 54 nsew signal input
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 wbs_adr_i[14]
port 55 nsew signal input
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 wbs_adr_i[15]
port 56 nsew signal input
flabel metal3 s 0 22176 800 22296 0 FreeSans 480 0 0 0 wbs_adr_i[16]
port 57 nsew signal input
flabel metal3 s 0 22992 800 23112 0 FreeSans 480 0 0 0 wbs_adr_i[17]
port 58 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 wbs_adr_i[18]
port 59 nsew signal input
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 wbs_adr_i[19]
port 60 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 wbs_adr_i[1]
port 61 nsew signal input
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 wbs_adr_i[20]
port 62 nsew signal input
flabel metal3 s 0 26256 800 26376 0 FreeSans 480 0 0 0 wbs_adr_i[21]
port 63 nsew signal input
flabel metal3 s 0 27072 800 27192 0 FreeSans 480 0 0 0 wbs_adr_i[22]
port 64 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 wbs_adr_i[23]
port 65 nsew signal input
flabel metal3 s 0 28704 800 28824 0 FreeSans 480 0 0 0 wbs_adr_i[24]
port 66 nsew signal input
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 wbs_adr_i[25]
port 67 nsew signal input
flabel metal3 s 0 30336 800 30456 0 FreeSans 480 0 0 0 wbs_adr_i[26]
port 68 nsew signal input
flabel metal3 s 0 31152 800 31272 0 FreeSans 480 0 0 0 wbs_adr_i[27]
port 69 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 wbs_adr_i[28]
port 70 nsew signal input
flabel metal3 s 0 32784 800 32904 0 FreeSans 480 0 0 0 wbs_adr_i[29]
port 71 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 wbs_adr_i[2]
port 72 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 wbs_adr_i[30]
port 73 nsew signal input
flabel metal3 s 0 34416 800 34536 0 FreeSans 480 0 0 0 wbs_adr_i[31]
port 74 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 wbs_adr_i[3]
port 75 nsew signal input
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 wbs_adr_i[4]
port 76 nsew signal input
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 wbs_adr_i[5]
port 77 nsew signal input
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 wbs_adr_i[6]
port 78 nsew signal input
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 wbs_adr_i[7]
port 79 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 wbs_adr_i[8]
port 80 nsew signal input
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 wbs_adr_i[9]
port 81 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 wbs_cyc_i
port 82 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 wbs_dat_i[0]
port 83 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 wbs_dat_i[10]
port 84 nsew signal input
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 wbs_dat_i[11]
port 85 nsew signal input
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 wbs_dat_i[12]
port 86 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 wbs_dat_i[13]
port 87 nsew signal input
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 wbs_dat_i[14]
port 88 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 wbs_dat_i[15]
port 89 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 wbs_dat_i[16]
port 90 nsew signal input
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 wbs_dat_i[17]
port 91 nsew signal input
flabel metal3 s 0 24216 800 24336 0 FreeSans 480 0 0 0 wbs_dat_i[18]
port 92 nsew signal input
flabel metal3 s 0 25032 800 25152 0 FreeSans 480 0 0 0 wbs_dat_i[19]
port 93 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 wbs_dat_i[1]
port 94 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 wbs_dat_i[20]
port 95 nsew signal input
flabel metal3 s 0 26664 800 26784 0 FreeSans 480 0 0 0 wbs_dat_i[21]
port 96 nsew signal input
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 wbs_dat_i[22]
port 97 nsew signal input
flabel metal3 s 0 28296 800 28416 0 FreeSans 480 0 0 0 wbs_dat_i[23]
port 98 nsew signal input
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 wbs_dat_i[24]
port 99 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 wbs_dat_i[25]
port 100 nsew signal input
flabel metal3 s 0 30744 800 30864 0 FreeSans 480 0 0 0 wbs_dat_i[26]
port 101 nsew signal input
flabel metal3 s 0 31560 800 31680 0 FreeSans 480 0 0 0 wbs_dat_i[27]
port 102 nsew signal input
flabel metal3 s 0 32376 800 32496 0 FreeSans 480 0 0 0 wbs_dat_i[28]
port 103 nsew signal input
flabel metal3 s 0 33192 800 33312 0 FreeSans 480 0 0 0 wbs_dat_i[29]
port 104 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 wbs_dat_i[2]
port 105 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 wbs_dat_i[30]
port 106 nsew signal input
flabel metal3 s 0 34824 800 34944 0 FreeSans 480 0 0 0 wbs_dat_i[31]
port 107 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 wbs_dat_i[3]
port 108 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 wbs_dat_i[4]
port 109 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 wbs_dat_i[5]
port 110 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 wbs_dat_i[6]
port 111 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 wbs_dat_i[7]
port 112 nsew signal input
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 wbs_dat_i[8]
port 113 nsew signal input
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 wbs_dat_i[9]
port 114 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 wbs_sel_i[0]
port 115 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 wbs_sel_i[1]
port 116 nsew signal input
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 wbs_sel_i[2]
port 117 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 wbs_sel_i[3]
port 118 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 wbs_stb_i
port 119 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 wbs_we_i
port 120 nsew signal input
flabel metal3 s 39200 5312 40000 5432 0 FreeSans 480 0 0 0 web0
port 121 nsew signal tristate
flabel metal3 s 39200 5992 40000 6112 0 FreeSans 480 0 0 0 wmask0[0]
port 122 nsew signal tristate
flabel metal3 s 39200 6672 40000 6792 0 FreeSans 480 0 0 0 wmask0[1]
port 123 nsew signal tristate
flabel metal3 s 39200 7352 40000 7472 0 FreeSans 480 0 0 0 wmask0[2]
port 124 nsew signal tristate
flabel metal3 s 39200 8032 40000 8152 0 FreeSans 480 0 0 0 wmask0[3]
port 125 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
