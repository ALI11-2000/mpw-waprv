magic
tech sky130B
magscale 1 2
timestamp 1661333512
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 2128 38824 37584
<< obsm2 >>
rect 1306 2139 38344 37573
<< metal3 >>
rect 39200 36592 40000 36712
rect 39200 35912 40000 36032
rect 39200 35232 40000 35352
rect 0 34824 800 34944
rect 0 34416 800 34536
rect 39200 34552 40000 34672
rect 0 34008 800 34128
rect 39200 33872 40000 33992
rect 0 33600 800 33720
rect 0 33192 800 33312
rect 39200 33192 40000 33312
rect 0 32784 800 32904
rect 0 32376 800 32496
rect 39200 32512 40000 32632
rect 0 31968 800 32088
rect 39200 31832 40000 31952
rect 0 31560 800 31680
rect 0 31152 800 31272
rect 39200 31152 40000 31272
rect 0 30744 800 30864
rect 0 30336 800 30456
rect 39200 30472 40000 30592
rect 0 29928 800 30048
rect 39200 29792 40000 29912
rect 0 29520 800 29640
rect 0 29112 800 29232
rect 39200 29112 40000 29232
rect 0 28704 800 28824
rect 0 28296 800 28416
rect 39200 28432 40000 28552
rect 0 27888 800 28008
rect 39200 27752 40000 27872
rect 0 27480 800 27600
rect 0 27072 800 27192
rect 39200 27072 40000 27192
rect 0 26664 800 26784
rect 0 26256 800 26376
rect 39200 26392 40000 26512
rect 0 25848 800 25968
rect 39200 25712 40000 25832
rect 0 25440 800 25560
rect 0 25032 800 25152
rect 39200 25032 40000 25152
rect 0 24624 800 24744
rect 0 24216 800 24336
rect 39200 24352 40000 24472
rect 0 23808 800 23928
rect 39200 23672 40000 23792
rect 0 23400 800 23520
rect 0 22992 800 23112
rect 39200 22992 40000 23112
rect 0 22584 800 22704
rect 0 22176 800 22296
rect 39200 22312 40000 22432
rect 0 21768 800 21888
rect 39200 21632 40000 21752
rect 0 21360 800 21480
rect 0 20952 800 21072
rect 39200 20952 40000 21072
rect 0 20544 800 20664
rect 0 20136 800 20256
rect 39200 20272 40000 20392
rect 0 19728 800 19848
rect 39200 19592 40000 19712
rect 0 19320 800 19440
rect 0 18912 800 19032
rect 39200 18912 40000 19032
rect 0 18504 800 18624
rect 0 18096 800 18216
rect 39200 18232 40000 18352
rect 0 17688 800 17808
rect 39200 17552 40000 17672
rect 0 17280 800 17400
rect 0 16872 800 16992
rect 39200 16872 40000 16992
rect 0 16464 800 16584
rect 0 16056 800 16176
rect 39200 16192 40000 16312
rect 0 15648 800 15768
rect 39200 15512 40000 15632
rect 0 15240 800 15360
rect 0 14832 800 14952
rect 39200 14832 40000 14952
rect 0 14424 800 14544
rect 0 14016 800 14136
rect 39200 14152 40000 14272
rect 0 13608 800 13728
rect 39200 13472 40000 13592
rect 0 13200 800 13320
rect 0 12792 800 12912
rect 39200 12792 40000 12912
rect 0 12384 800 12504
rect 0 11976 800 12096
rect 39200 12112 40000 12232
rect 0 11568 800 11688
rect 39200 11432 40000 11552
rect 0 11160 800 11280
rect 0 10752 800 10872
rect 39200 10752 40000 10872
rect 0 10344 800 10464
rect 0 9936 800 10056
rect 39200 10072 40000 10192
rect 0 9528 800 9648
rect 39200 9392 40000 9512
rect 0 9120 800 9240
rect 0 8712 800 8832
rect 39200 8712 40000 8832
rect 0 8304 800 8424
rect 0 7896 800 8016
rect 39200 8032 40000 8152
rect 0 7488 800 7608
rect 39200 7352 40000 7472
rect 0 7080 800 7200
rect 0 6672 800 6792
rect 39200 6672 40000 6792
rect 0 6264 800 6384
rect 0 5856 800 5976
rect 39200 5992 40000 6112
rect 0 5448 800 5568
rect 39200 5312 40000 5432
rect 0 5040 800 5160
rect 39200 4632 40000 4752
rect 39200 3952 40000 4072
rect 39200 3272 40000 3392
<< obsm3 >>
rect 800 36792 39200 37569
rect 800 36512 39120 36792
rect 800 36112 39200 36512
rect 800 35832 39120 36112
rect 800 35432 39200 35832
rect 800 35152 39120 35432
rect 800 35024 39200 35152
rect 880 34752 39200 35024
rect 880 34744 39120 34752
rect 800 34616 39120 34744
rect 880 34472 39120 34616
rect 880 34336 39200 34472
rect 800 34208 39200 34336
rect 880 34072 39200 34208
rect 880 33928 39120 34072
rect 800 33800 39120 33928
rect 880 33792 39120 33800
rect 880 33520 39200 33792
rect 800 33392 39200 33520
rect 880 33112 39120 33392
rect 800 32984 39200 33112
rect 880 32712 39200 32984
rect 880 32704 39120 32712
rect 800 32576 39120 32704
rect 880 32432 39120 32576
rect 880 32296 39200 32432
rect 800 32168 39200 32296
rect 880 32032 39200 32168
rect 880 31888 39120 32032
rect 800 31760 39120 31888
rect 880 31752 39120 31760
rect 880 31480 39200 31752
rect 800 31352 39200 31480
rect 880 31072 39120 31352
rect 800 30944 39200 31072
rect 880 30672 39200 30944
rect 880 30664 39120 30672
rect 800 30536 39120 30664
rect 880 30392 39120 30536
rect 880 30256 39200 30392
rect 800 30128 39200 30256
rect 880 29992 39200 30128
rect 880 29848 39120 29992
rect 800 29720 39120 29848
rect 880 29712 39120 29720
rect 880 29440 39200 29712
rect 800 29312 39200 29440
rect 880 29032 39120 29312
rect 800 28904 39200 29032
rect 880 28632 39200 28904
rect 880 28624 39120 28632
rect 800 28496 39120 28624
rect 880 28352 39120 28496
rect 880 28216 39200 28352
rect 800 28088 39200 28216
rect 880 27952 39200 28088
rect 880 27808 39120 27952
rect 800 27680 39120 27808
rect 880 27672 39120 27680
rect 880 27400 39200 27672
rect 800 27272 39200 27400
rect 880 26992 39120 27272
rect 800 26864 39200 26992
rect 880 26592 39200 26864
rect 880 26584 39120 26592
rect 800 26456 39120 26584
rect 880 26312 39120 26456
rect 880 26176 39200 26312
rect 800 26048 39200 26176
rect 880 25912 39200 26048
rect 880 25768 39120 25912
rect 800 25640 39120 25768
rect 880 25632 39120 25640
rect 880 25360 39200 25632
rect 800 25232 39200 25360
rect 880 24952 39120 25232
rect 800 24824 39200 24952
rect 880 24552 39200 24824
rect 880 24544 39120 24552
rect 800 24416 39120 24544
rect 880 24272 39120 24416
rect 880 24136 39200 24272
rect 800 24008 39200 24136
rect 880 23872 39200 24008
rect 880 23728 39120 23872
rect 800 23600 39120 23728
rect 880 23592 39120 23600
rect 880 23320 39200 23592
rect 800 23192 39200 23320
rect 880 22912 39120 23192
rect 800 22784 39200 22912
rect 880 22512 39200 22784
rect 880 22504 39120 22512
rect 800 22376 39120 22504
rect 880 22232 39120 22376
rect 880 22096 39200 22232
rect 800 21968 39200 22096
rect 880 21832 39200 21968
rect 880 21688 39120 21832
rect 800 21560 39120 21688
rect 880 21552 39120 21560
rect 880 21280 39200 21552
rect 800 21152 39200 21280
rect 880 20872 39120 21152
rect 800 20744 39200 20872
rect 880 20472 39200 20744
rect 880 20464 39120 20472
rect 800 20336 39120 20464
rect 880 20192 39120 20336
rect 880 20056 39200 20192
rect 800 19928 39200 20056
rect 880 19792 39200 19928
rect 880 19648 39120 19792
rect 800 19520 39120 19648
rect 880 19512 39120 19520
rect 880 19240 39200 19512
rect 800 19112 39200 19240
rect 880 18832 39120 19112
rect 800 18704 39200 18832
rect 880 18432 39200 18704
rect 880 18424 39120 18432
rect 800 18296 39120 18424
rect 880 18152 39120 18296
rect 880 18016 39200 18152
rect 800 17888 39200 18016
rect 880 17752 39200 17888
rect 880 17608 39120 17752
rect 800 17480 39120 17608
rect 880 17472 39120 17480
rect 880 17200 39200 17472
rect 800 17072 39200 17200
rect 880 16792 39120 17072
rect 800 16664 39200 16792
rect 880 16392 39200 16664
rect 880 16384 39120 16392
rect 800 16256 39120 16384
rect 880 16112 39120 16256
rect 880 15976 39200 16112
rect 800 15848 39200 15976
rect 880 15712 39200 15848
rect 880 15568 39120 15712
rect 800 15440 39120 15568
rect 880 15432 39120 15440
rect 880 15160 39200 15432
rect 800 15032 39200 15160
rect 880 14752 39120 15032
rect 800 14624 39200 14752
rect 880 14352 39200 14624
rect 880 14344 39120 14352
rect 800 14216 39120 14344
rect 880 14072 39120 14216
rect 880 13936 39200 14072
rect 800 13808 39200 13936
rect 880 13672 39200 13808
rect 880 13528 39120 13672
rect 800 13400 39120 13528
rect 880 13392 39120 13400
rect 880 13120 39200 13392
rect 800 12992 39200 13120
rect 880 12712 39120 12992
rect 800 12584 39200 12712
rect 880 12312 39200 12584
rect 880 12304 39120 12312
rect 800 12176 39120 12304
rect 880 12032 39120 12176
rect 880 11896 39200 12032
rect 800 11768 39200 11896
rect 880 11632 39200 11768
rect 880 11488 39120 11632
rect 800 11360 39120 11488
rect 880 11352 39120 11360
rect 880 11080 39200 11352
rect 800 10952 39200 11080
rect 880 10672 39120 10952
rect 800 10544 39200 10672
rect 880 10272 39200 10544
rect 880 10264 39120 10272
rect 800 10136 39120 10264
rect 880 9992 39120 10136
rect 880 9856 39200 9992
rect 800 9728 39200 9856
rect 880 9592 39200 9728
rect 880 9448 39120 9592
rect 800 9320 39120 9448
rect 880 9312 39120 9320
rect 880 9040 39200 9312
rect 800 8912 39200 9040
rect 880 8632 39120 8912
rect 800 8504 39200 8632
rect 880 8232 39200 8504
rect 880 8224 39120 8232
rect 800 8096 39120 8224
rect 880 7952 39120 8096
rect 880 7816 39200 7952
rect 800 7688 39200 7816
rect 880 7552 39200 7688
rect 880 7408 39120 7552
rect 800 7280 39120 7408
rect 880 7272 39120 7280
rect 880 7000 39200 7272
rect 800 6872 39200 7000
rect 880 6592 39120 6872
rect 800 6464 39200 6592
rect 880 6192 39200 6464
rect 880 6184 39120 6192
rect 800 6056 39120 6184
rect 880 5912 39120 6056
rect 880 5776 39200 5912
rect 800 5648 39200 5776
rect 880 5512 39200 5648
rect 880 5368 39120 5512
rect 800 5240 39120 5368
rect 880 5232 39120 5240
rect 880 4960 39200 5232
rect 800 4832 39200 4960
rect 800 4552 39120 4832
rect 800 4152 39200 4552
rect 800 3872 39120 4152
rect 800 3472 39200 3872
rect 800 3192 39120 3472
rect 800 2143 39200 3192
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 2635 24107 2701 27709
<< labels >>
rlabel metal3 s 39200 30472 40000 30592 6 addr0[0]
port 1 nsew signal output
rlabel metal3 s 39200 31152 40000 31272 6 addr0[1]
port 2 nsew signal output
rlabel metal3 s 39200 31832 40000 31952 6 addr0[2]
port 3 nsew signal output
rlabel metal3 s 39200 32512 40000 32632 6 addr0[3]
port 4 nsew signal output
rlabel metal3 s 39200 33192 40000 33312 6 addr0[4]
port 5 nsew signal output
rlabel metal3 s 39200 33872 40000 33992 6 addr0[5]
port 6 nsew signal output
rlabel metal3 s 39200 34552 40000 34672 6 addr0[6]
port 7 nsew signal output
rlabel metal3 s 39200 35232 40000 35352 6 addr0[7]
port 8 nsew signal output
rlabel metal3 s 39200 35912 40000 36032 6 addr0[8]
port 9 nsew signal output
rlabel metal3 s 39200 3952 40000 4072 6 clk0
port 10 nsew signal output
rlabel metal3 s 39200 4632 40000 4752 6 csb0
port 11 nsew signal output
rlabel metal3 s 39200 8712 40000 8832 6 din0[0]
port 12 nsew signal output
rlabel metal3 s 39200 15512 40000 15632 6 din0[10]
port 13 nsew signal output
rlabel metal3 s 39200 16192 40000 16312 6 din0[11]
port 14 nsew signal output
rlabel metal3 s 39200 16872 40000 16992 6 din0[12]
port 15 nsew signal output
rlabel metal3 s 39200 17552 40000 17672 6 din0[13]
port 16 nsew signal output
rlabel metal3 s 39200 18232 40000 18352 6 din0[14]
port 17 nsew signal output
rlabel metal3 s 39200 18912 40000 19032 6 din0[15]
port 18 nsew signal output
rlabel metal3 s 39200 19592 40000 19712 6 din0[16]
port 19 nsew signal output
rlabel metal3 s 39200 20272 40000 20392 6 din0[17]
port 20 nsew signal output
rlabel metal3 s 39200 20952 40000 21072 6 din0[18]
port 21 nsew signal output
rlabel metal3 s 39200 21632 40000 21752 6 din0[19]
port 22 nsew signal output
rlabel metal3 s 39200 9392 40000 9512 6 din0[1]
port 23 nsew signal output
rlabel metal3 s 39200 22312 40000 22432 6 din0[20]
port 24 nsew signal output
rlabel metal3 s 39200 22992 40000 23112 6 din0[21]
port 25 nsew signal output
rlabel metal3 s 39200 23672 40000 23792 6 din0[22]
port 26 nsew signal output
rlabel metal3 s 39200 24352 40000 24472 6 din0[23]
port 27 nsew signal output
rlabel metal3 s 39200 25032 40000 25152 6 din0[24]
port 28 nsew signal output
rlabel metal3 s 39200 25712 40000 25832 6 din0[25]
port 29 nsew signal output
rlabel metal3 s 39200 26392 40000 26512 6 din0[26]
port 30 nsew signal output
rlabel metal3 s 39200 27072 40000 27192 6 din0[27]
port 31 nsew signal output
rlabel metal3 s 39200 27752 40000 27872 6 din0[28]
port 32 nsew signal output
rlabel metal3 s 39200 28432 40000 28552 6 din0[29]
port 33 nsew signal output
rlabel metal3 s 39200 10072 40000 10192 6 din0[2]
port 34 nsew signal output
rlabel metal3 s 39200 29112 40000 29232 6 din0[30]
port 35 nsew signal output
rlabel metal3 s 39200 29792 40000 29912 6 din0[31]
port 36 nsew signal output
rlabel metal3 s 39200 10752 40000 10872 6 din0[3]
port 37 nsew signal output
rlabel metal3 s 39200 11432 40000 11552 6 din0[4]
port 38 nsew signal output
rlabel metal3 s 39200 12112 40000 12232 6 din0[5]
port 39 nsew signal output
rlabel metal3 s 39200 12792 40000 12912 6 din0[6]
port 40 nsew signal output
rlabel metal3 s 39200 13472 40000 13592 6 din0[7]
port 41 nsew signal output
rlabel metal3 s 39200 14152 40000 14272 6 din0[8]
port 42 nsew signal output
rlabel metal3 s 39200 14832 40000 14952 6 din0[9]
port 43 nsew signal output
rlabel metal3 s 39200 3272 40000 3392 6 imem_rd_cs1
port 44 nsew signal output
rlabel metal3 s 39200 36592 40000 36712 6 processor_reset
port 45 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 46 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 46 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 47 nsew ground bidirectional
rlabel metal3 s 0 5040 800 5160 6 wb_clk_i
port 48 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 wb_rst_i
port 49 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 wbs_ack_o
port 50 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 wbs_adr_i[0]
port 51 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 wbs_adr_i[10]
port 52 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wbs_adr_i[11]
port 53 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 wbs_adr_i[12]
port 54 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 wbs_adr_i[13]
port 55 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 wbs_adr_i[14]
port 56 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 wbs_adr_i[15]
port 57 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 wbs_adr_i[16]
port 58 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 wbs_adr_i[17]
port 59 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_adr_i[18]
port 60 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 wbs_adr_i[19]
port 61 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 wbs_adr_i[1]
port 62 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 wbs_adr_i[20]
port 63 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 wbs_adr_i[21]
port 64 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 wbs_adr_i[22]
port 65 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 wbs_adr_i[23]
port 66 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 wbs_adr_i[24]
port 67 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 wbs_adr_i[25]
port 68 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wbs_adr_i[26]
port 69 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 wbs_adr_i[27]
port 70 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 wbs_adr_i[28]
port 71 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 wbs_adr_i[29]
port 72 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 wbs_adr_i[2]
port 73 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 wbs_adr_i[30]
port 74 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 wbs_adr_i[31]
port 75 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 wbs_adr_i[3]
port 76 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 wbs_adr_i[4]
port 77 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 wbs_adr_i[5]
port 78 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 wbs_adr_i[6]
port 79 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 wbs_adr_i[7]
port 80 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wbs_adr_i[8]
port 81 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wbs_adr_i[9]
port 82 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 wbs_cyc_i
port 83 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 wbs_dat_i[0]
port 84 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wbs_dat_i[10]
port 85 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 wbs_dat_i[11]
port 86 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 wbs_dat_i[12]
port 87 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 wbs_dat_i[13]
port 88 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 wbs_dat_i[14]
port 89 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_i[15]
port 90 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 wbs_dat_i[16]
port 91 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 wbs_dat_i[17]
port 92 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 wbs_dat_i[18]
port 93 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 wbs_dat_i[19]
port 94 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 wbs_dat_i[1]
port 95 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_dat_i[20]
port 96 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 wbs_dat_i[21]
port 97 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wbs_dat_i[22]
port 98 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 wbs_dat_i[23]
port 99 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wbs_dat_i[24]
port 100 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 wbs_dat_i[25]
port 101 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wbs_dat_i[26]
port 102 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wbs_dat_i[27]
port 103 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 wbs_dat_i[28]
port 104 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 wbs_dat_i[29]
port 105 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 wbs_dat_i[2]
port 106 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 wbs_dat_i[30]
port 107 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 wbs_dat_i[31]
port 108 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_dat_i[3]
port 109 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 wbs_dat_i[4]
port 110 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 wbs_dat_i[5]
port 111 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 wbs_dat_i[6]
port 112 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 wbs_dat_i[7]
port 113 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 wbs_dat_i[8]
port 114 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wbs_dat_i[9]
port 115 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 wbs_sel_i[0]
port 116 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wbs_sel_i[1]
port 117 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 wbs_sel_i[2]
port 118 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 wbs_sel_i[3]
port 119 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 wbs_stb_i
port 120 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 wbs_we_i
port 121 nsew signal input
rlabel metal3 s 39200 5312 40000 5432 6 web0
port 122 nsew signal output
rlabel metal3 s 39200 5992 40000 6112 6 wmask0[0]
port 123 nsew signal output
rlabel metal3 s 39200 6672 40000 6792 6 wmask0[1]
port 124 nsew signal output
rlabel metal3 s 39200 7352 40000 7472 6 wmask0[2]
port 125 nsew signal output
rlabel metal3 s 39200 8032 40000 8152 6 wmask0[3]
port 126 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 873536
string GDS_FILE /home/ali11-2000/efabless/mpw-waprv/openlane/wb_interface/runs/22_08_24_14_30/results/signoff/wb_interface.magic.gds
string GDS_START 107132
<< end >>

